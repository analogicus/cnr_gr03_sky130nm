*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TOPLEVEL_lpe.spi
.include ../../../work/lpe/M3_lpe.spi
#else
.include ../../../work/xsch/TOPLEVEL.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

*.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0 dc 0
VDD  VDD_1V8  VSS  dc 1.8
Vclk clk VSS PULSE(0 1.8 0.0 2NS 2NS 12.5NS 25NS)
*VRST VRST VSS PULSE(0 1.8 0.0 2NS 2NS 10US 50US)
*IBIAS VDD IBIAS dc 2u

*VRST VRST VSS dc 0
Vtest rst VSS dc 0

    
*-----------------------------------------------------------------
* DUT xschem
*-----------------------------------------------------------------
*.subckt TOPLEVEL VDD VSS VOUT VRST
XDUT VDD_1V8 VSS VOUT rst2 TOPLEVEL
adut [clk VOUT rst] [rst2 d7 d6 d5 d4 d3 d2 d1 d0]  null dut
.model dut d_cosim simulation="../dtt.so"


*-----------------------------------------------------------------
* DUT lay
*-----------------------------------------------------------------
*.subckt M3 clk data_out[5] in data_out[0] data_out[2] data_out[7] data_out[4] data_out[6] data_out[1] rst data_out[3] rst_cap VPWR VGND
*xadut clk d5 VOUT d0 d2 d7 d4 d6 d1 rst2 d3 rst VDD VSS M3



*R11 rst2 rst 10k
R10 rst2 VSS 1M

R1 d1 VSS 1M
R2 d2 VSS 1M
R3 d3 VSS 1M
R4 d4 VSS 1M
R5 d5 VSS 1M
R6 d6 VSS 1M
R7 d7 VSS 1M
R0 d0 VSS 1M



*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

*.save all

*TOPLEVEL valuescat
.save v(VOUT) v(VRST) v(XDUT.VREF) v(XDUT.I_PTAT) 

*Milestone 1 values
.save v(XDUT.X1.OTA_OUT) v(XDUT.X1.VD1) v(XDUT.X1.VR1)

.save v(d0) v(d1) v(d2) v(d3) v(d4) v(d5) v(d6) v(d7)
.save v(clk) v(rst2)
*.save all

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

*save @m.xdut.x3.x7.xm1.msky130_fd_pr__pfet_01v8[id]


optran 0 0 0 10n 10u 0 


option TEMP=27
tran 10000m 475u 400u 100u
write {cicname}_27.raw


exit

.endc

.end
