magic
tech sky130B
magscale 1 2
timestamp 1712309541
<< locali >>
rect 422 4960 622 5346
rect 422 4760 18469 4960
rect 18669 4760 30184 4960
rect 27332 4400 29546 4600
rect 29346 3726 29546 4400
rect 30346 3726 30546 4160
rect 29346 3526 30558 3726
<< metal2 >>
rect 26258 17502 26322 17708
rect 26253 17446 26262 17502
rect 26318 17446 26327 17502
rect 26258 17442 26322 17446
rect 28894 13988 28958 14226
rect 28894 13915 28958 13924
rect 7264 8704 7328 8713
rect 7264 8631 7328 8640
rect 27036 8474 27356 8510
rect 27328 6352 27392 6361
rect 22268 6288 27328 6352
rect 27392 6288 28594 6352
rect 28658 6288 28664 6352
rect 27328 6279 27392 6288
rect 7582 5150 7642 5159
rect 7582 5081 7642 5090
<< via2 >>
rect 26262 17446 26318 17502
rect 28894 13924 28958 13988
rect 7264 8640 7328 8704
rect 27328 6288 27392 6352
rect 7582 5090 7642 5150
<< metal3 >>
rect 26257 17506 26323 17507
rect 26200 17502 26490 17506
rect 26200 17446 26262 17502
rect 26318 17446 26490 17502
rect 26200 17442 26490 17446
rect 26257 17441 26323 17442
rect 28889 13988 28963 13993
rect 26118 13924 28894 13988
rect 28958 13924 28963 13988
rect 26158 8872 26219 13924
rect 28889 13919 28963 13924
rect 7259 8704 7333 8709
rect 7259 8640 7264 8704
rect 7328 8640 7333 8704
rect 7259 8635 7333 8640
rect 7264 8548 7328 8635
rect 7258 8484 7264 8548
rect 7328 8484 7334 8548
rect 7580 5356 7644 5362
rect 26158 5356 26218 8872
rect 27323 6352 27397 6357
rect 27323 6288 27328 6352
rect 27392 6288 27397 6352
rect 27323 6283 27397 6288
rect 27328 5786 27392 6283
rect 26150 5292 26156 5356
rect 26220 5292 26226 5356
rect 7580 5286 7644 5292
rect 7582 5155 7642 5286
rect 7577 5150 7647 5155
rect 7577 5090 7582 5150
rect 7642 5090 7647 5150
rect 7577 5085 7647 5090
<< via3 >>
rect 7264 8484 7328 8548
rect 7580 5292 7644 5356
rect 26156 5292 26220 5356
<< metal4 >>
rect 7263 8548 7329 8549
rect 7263 8484 7264 8548
rect 7328 8484 27510 8548
rect 7263 8483 7329 8484
rect 7579 5356 7645 5357
rect 7579 5292 7580 5356
rect 7644 5354 7645 5356
rect 26155 5356 26221 5357
rect 26155 5354 26156 5356
rect 7644 5294 26156 5354
rect 7644 5292 7645 5294
rect 7579 5291 7645 5292
rect 26155 5292 26156 5294
rect 26220 5292 26221 5356
rect 26155 5291 26221 5292
use MILESTONE1  MILESTONE1_0
timestamp 1712303455
transform 1 0 -12348 0 1 4600
box 12340 -4600 39920 6836
use MILESTONE2  MILESTONE2_0
timestamp 1712303529
transform 0 -1 30538 1 0 5654
box -5400 -11400 18492 7028
<< labels >>
flabel metal2 27036 8474 27356 8510 0 FreeSans 800 0 0 0 VRST
port 4 nsew
flabel locali 29346 3526 29546 4600 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel metal2 26258 17502 26322 17708 0 FreeSans 800 0 0 0 VOUT
port 3 nsew
flabel locali 422 4760 622 5346 0 FreeSans 800 0 0 0 VSS
port 2 nsew
flabel metal3 27328 5786 27392 6288 0 FreeSans 1600 0 0 0 IBIAS
port 7 nsew
<< end >>
