*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/BIAS_lpe.spi
#else
.include ../../../work/xsch/BIAS.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0 dc 0
VDD  VDD_1V8  VSS  dc 1.8
V1 IBIAS1 VSS dc 0
V2 IBIAS2 VSS dc 0

*-----------------------------------------------------------------
* DUT

XDUT VDD_1V8 VSS IBIAS1 IBIAS2 BIAS

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save i(V0)
#else
.save i(v1) v(VDD_1V8) v(VSS) i(v2)
*.save all
#endif


*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

save @m.xdut.x7.xm1.msky130_fd_pr__pfet_01v8[id]

optran 0 0 0 100n 10u 0

#ifdef Debug
tran 10p 1n 1p
*quit
#else
tran 10m 10m 400u
write
quit
#endif

.endc

.end
