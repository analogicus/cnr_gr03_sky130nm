magic
tech sky130B
magscale 1 2
timestamp 1712845386
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 5144 -1 0 1256
box -184 -124 1336 2168
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 1604 0 1 1024
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_1
timestamp 1695852000
transform 1 0 1604 0 1 3064
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_2
timestamp 1695852000
transform 1 0 1604 0 1 2044
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_3
timestamp 1695852000
transform 1 0 -36 0 1 4
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_4
timestamp 1695852000
transform 1 0 -36 0 1 3064
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_5
timestamp 1695852000
transform 1 0 -36 0 1 2044
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_6
timestamp 1695852000
transform 1 0 -36 0 1 1024
box -184 -124 1528 1016
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 3324 0 1 4
box -184 -124 1528 1016
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_1
timestamp 1695852000
transform 1 0 3324 0 1 3064
box -184 -124 1528 1016
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_2
timestamp 1695852000
transform 1 0 3324 0 1 2044
box -184 -124 1528 1016
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_3
timestamp 1695852000
transform 1 0 3324 0 1 1024
box -184 -124 1528 1016
use CNRATR_PCH_12C1F2  CNRATR_PCH_12C1F2_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 5884 -1 0 3796
box -184 -124 2296 613
use CNRATR_PCH_12C1F2  CNRATR_PCH_12C1F2_1
timestamp 1695852000
transform 0 1 5264 -1 0 3796
box -184 -124 2296 613
use SUNTR_RPPO8  SUNTR_RPPO8_0 ~/aicex/ip/cnr_gr03_sky130nm/design/SUN_TR_SKY130NM
timestamp 1712819652
transform 1 0 -5540 0 1 -60
box 0 0 5264 4236
<< end >>
