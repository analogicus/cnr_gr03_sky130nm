magic
tech sky130B
magscale 1 2
timestamp 1711370500
<< locali >>
rect 13111 4512 15356 4584
rect 16211 4512 18456 4584
rect 12708 3697 12863 3783
rect 18697 3697 18849 3783
rect 19437 3697 19585 3783
rect 12708 3154 12794 3697
rect 13052 3440 15792 3497
rect 15850 3440 18488 3497
rect 18763 3183 18849 3697
rect 19069 3432 19071 3491
rect 19131 3432 19204 3491
rect 13157 3102 18374 3183
rect 13157 3097 16268 3102
rect 16332 3097 18374 3102
rect 18763 3097 19103 3183
rect 19499 3154 19585 3697
rect 14171 2152 14536 2224
rect 14791 2152 15176 2224
rect 15429 2222 15857 2224
rect 15186 2150 15857 2222
rect 16051 2144 16476 2216
rect 36279 1904 36351 2376
rect 37567 1899 37639 2376
rect 16677 1357 16835 1443
rect 14112 1080 15272 1136
rect 15328 1080 15612 1136
rect 15668 1080 16528 1136
rect 14243 737 14483 823
rect 14863 737 15123 823
rect 15503 806 15763 823
rect 15503 754 15614 806
rect 15666 754 15763 806
rect 15503 737 15763 754
rect 16123 737 16383 823
rect 16749 794 16835 1357
rect 17891 360 17990 985
rect 18045 884 18117 1121
rect 35226 360 35325 945
rect 37711 846 37965 945
rect 38029 844 38101 1081
rect 14100 290 39896 360
rect 14100 257 19230 290
rect 13749 199 19230 257
rect 13749 -406 13807 199
rect 14100 190 19230 199
rect 19330 190 22110 290
rect 22210 270 39896 290
rect 22210 190 31050 270
rect 14100 170 31050 190
rect 31150 170 39896 270
rect 14100 160 39896 170
rect 17891 151 17990 160
rect 14100 -74 19500 0
rect 14100 -126 15614 -74
rect 15666 -126 16274 -74
rect 16326 -126 19500 -74
rect 14100 -200 19500 -126
rect 34400 -200 39880 0
rect 13419 -641 13491 -424
rect 13596 -464 13809 -406
rect 19044 -492 19224 -380
rect 19336 -492 19536 -380
rect 21944 -492 22104 -380
rect 22216 -492 22436 -380
rect 30892 -492 31044 -380
rect 31156 -492 31356 -380
rect 22056 -961 22064 -880
rect 14779 -1516 15256 -1444
rect 31805 -1497 32036 -1442
rect 31915 -1607 32036 -1497
rect 31805 -1662 32036 -1607
rect 14779 -1921 15276 -1849
<< viali >>
rect 12973 4040 13024 4104
rect 13580 4053 13620 4093
rect 14200 4053 14240 4093
rect 14840 4053 14880 4093
rect 15460 4053 15500 4093
rect 16060 4040 16124 4104
rect 16674 4046 16726 4098
rect 17294 4046 17346 4098
rect 17914 4046 17966 4098
rect 18534 4046 18586 4098
rect 19270 4040 19334 4104
rect 15792 3440 15850 3497
rect 19071 3432 19131 3491
rect 16268 3038 16332 3102
rect 14032 1680 14084 1744
rect 14665 1680 14704 1744
rect 15272 1680 15310 1744
rect 15892 1680 15956 1744
rect 16518 1680 16561 1744
rect 34234 1688 34298 1752
rect 15612 1080 15668 1136
rect 15614 754 15666 806
rect 25070 1272 25134 1336
rect 26670 1272 26734 1336
rect 19230 190 19330 290
rect 22110 190 22210 290
rect 31050 170 31150 270
rect 15614 -126 15666 -74
rect 16274 -126 16326 -74
rect 19224 -492 19336 -380
rect 22104 -492 22216 -380
rect 31044 -492 31156 -380
rect 17253 -1067 17307 -1013
rect 18254 -1086 18306 -1034
rect 20123 -1057 20157 -1023
rect 21299 -1162 21456 -942
rect 22927 -1124 23072 -979
rect 30258 -1162 30404 -942
rect 31873 -1119 32007 -985
rect 39113 -1067 39167 -1013
<< metal1 >>
rect 12967 4110 13030 4116
rect 16054 4110 16130 4116
rect 19264 4110 19340 4116
rect 12967 4104 12978 4110
rect 12967 4040 12973 4104
rect 12967 4034 12978 4040
rect 13030 4034 13036 4110
rect 13574 4099 13626 4105
rect 13574 4041 13626 4047
rect 14194 4099 14246 4105
rect 14194 4041 14246 4047
rect 14834 4099 14886 4105
rect 15454 4099 15506 4105
rect 15129 4047 15135 4099
rect 15187 4047 15193 4099
rect 14834 4041 14886 4047
rect 12967 4028 13030 4034
rect 15142 2933 15181 4047
rect 15454 4041 15506 4047
rect 16054 4104 16066 4110
rect 16054 4040 16060 4104
rect 16054 4034 16066 4040
rect 16130 4034 16136 4110
rect 16668 4104 16732 4110
rect 17288 4104 17352 4110
rect 17042 4040 17048 4104
rect 17112 4040 17118 4104
rect 16668 4034 16732 4040
rect 16054 4028 16130 4034
rect 15780 3497 15862 3503
rect 15780 3491 15792 3497
rect 15850 3491 15862 3497
rect 15780 3434 15786 3491
rect 15856 3434 15862 3491
rect 15786 3428 15856 3434
rect 16256 3102 16344 3108
rect 16256 3038 16268 3102
rect 16332 3038 16344 3102
rect 16256 3032 16344 3038
rect 15136 2927 15188 2933
rect 15136 2869 15188 2875
rect 14026 1750 14090 1756
rect 14659 1750 14710 1756
rect 15266 1750 15316 1756
rect 15886 1750 15962 1756
rect 14026 1744 14038 1750
rect 14026 1680 14032 1744
rect 14026 1674 14038 1680
rect 14090 1674 14096 1750
rect 14653 1674 14659 1750
rect 14711 1674 14717 1750
rect 14948 1686 14954 1738
rect 15006 1686 15012 1738
rect 14026 1668 14090 1674
rect 14659 1668 14710 1674
rect 14954 546 15006 1686
rect 15259 1674 15265 1750
rect 15317 1674 15323 1750
rect 15880 1674 15886 1750
rect 15938 1744 15962 1750
rect 15956 1680 15962 1744
rect 15938 1674 15962 1680
rect 15266 1668 15316 1674
rect 15886 1668 15962 1674
rect 15606 1142 15674 1148
rect 15600 1086 15606 1142
rect 15674 1086 15680 1142
rect 15600 1080 15612 1086
rect 15668 1080 15680 1086
rect 15600 1074 15680 1080
rect 15608 806 15672 818
rect 15608 754 15614 806
rect 15666 754 15672 806
rect 14948 494 14954 546
rect 15006 494 15012 546
rect 15608 -74 15672 754
rect 16268 -68 16332 3032
rect 17048 2292 17112 4040
rect 17288 4034 17352 4040
rect 17908 4104 17972 4110
rect 17908 4034 17972 4040
rect 18528 4104 18592 4110
rect 18528 4034 18592 4040
rect 19264 4104 19276 4110
rect 19264 4040 19270 4104
rect 19264 4034 19276 4040
rect 19340 4034 19346 4110
rect 19264 4028 19340 4034
rect 19059 3491 19143 3497
rect 19059 3485 19071 3491
rect 19131 3485 19143 3491
rect 19059 3426 19065 3485
rect 19137 3426 19143 3485
rect 19065 3420 19137 3426
rect 17414 2931 17466 2934
rect 16512 1750 16567 1756
rect 16506 1674 16512 1750
rect 16564 1674 16570 1750
rect 16512 1668 16567 1674
rect 15608 -126 15614 -74
rect 15666 -126 15672 -74
rect 15608 -138 15672 -126
rect 16262 -74 16338 -68
rect 16262 -126 16274 -74
rect 16326 -126 16338 -74
rect 16262 -132 16338 -126
rect 17048 -268 17112 2228
rect 17409 2928 17471 2931
rect 17409 2876 17414 2928
rect 17466 2876 17471 2928
rect 17409 2118 17471 2876
rect 36030 2567 36096 2579
rect 36030 2501 36951 2567
rect 17409 2112 17472 2118
rect 17409 2043 17472 2049
rect 17409 1693 17471 2043
rect 34228 1758 34304 1764
rect 34228 1752 34240 1758
rect 17407 1553 17473 1693
rect 34228 1688 34234 1752
rect 34228 1682 34240 1688
rect 34304 1682 34310 1758
rect 36030 1751 36096 2501
rect 36885 1751 36951 2501
rect 36030 1685 36951 1751
rect 34228 1676 34304 1682
rect 17401 1487 17407 1553
rect 17473 1487 17479 1553
rect 18480 1487 18486 1553
rect 18552 1487 18558 1553
rect 37127 1513 37193 1519
rect 37118 1447 37127 1493
rect 37118 1441 37193 1447
rect 25064 1342 25140 1348
rect 26664 1342 26740 1348
rect 25058 1266 25064 1342
rect 25128 1336 25140 1342
rect 25134 1272 25140 1336
rect 25128 1266 25140 1272
rect 26658 1278 26664 1342
rect 26740 1278 26746 1342
rect 26658 1272 26670 1278
rect 26734 1272 26746 1278
rect 26658 1266 26746 1272
rect 25064 1260 25140 1266
rect 37118 593 37184 1441
rect 37327 1407 38436 1473
rect 20108 494 20114 546
rect 20166 494 20172 546
rect 37118 521 37184 527
rect 39107 593 39173 599
rect 19224 290 19336 302
rect 19224 190 19230 290
rect 19330 190 19336 290
rect 17042 -332 17048 -268
rect 17112 -332 17118 -268
rect 18242 -332 18248 -268
rect 18312 -332 18318 -268
rect 13147 -1113 14196 -1047
rect 15612 -1073 15618 -1007
rect 15684 -1073 15690 -1007
rect 17241 -1073 17247 -1007
rect 17313 -1073 17319 -1007
rect 18248 -1034 18312 -332
rect 19224 -374 19336 190
rect 19212 -380 19348 -374
rect 19212 -492 19224 -380
rect 19336 -492 19348 -380
rect 19212 -498 19348 -492
rect 20120 -1011 20160 494
rect 22104 290 22216 302
rect 22104 190 22110 290
rect 22210 190 22216 290
rect 22104 -374 22216 190
rect 31038 270 31162 276
rect 31038 170 31050 270
rect 31150 170 31162 270
rect 31038 164 31162 170
rect 31044 -374 31156 164
rect 22092 -380 22228 -374
rect 22092 -492 22104 -380
rect 22216 -492 22228 -380
rect 22092 -498 22228 -492
rect 31032 -380 31168 -374
rect 31032 -492 31044 -380
rect 31156 -492 31168 -380
rect 31032 -498 31168 -492
rect 21293 -936 21462 -930
rect 30252 -936 30410 -930
rect 21293 -942 21305 -936
rect 18248 -1086 18254 -1034
rect 18306 -1086 18312 -1034
rect 20117 -1023 20163 -1011
rect 20117 -1057 20123 -1023
rect 20157 -1057 20163 -1023
rect 20117 -1069 20163 -1057
rect 18248 -1098 18312 -1086
rect 21293 -1162 21299 -942
rect 21293 -1168 21305 -1162
rect 21462 -1168 21468 -936
rect 30252 -942 30264 -936
rect 22921 -973 23078 -967
rect 22921 -1136 23078 -1130
rect 30252 -1162 30258 -942
rect 30252 -1168 30264 -1162
rect 30410 -1168 30416 -936
rect 31867 -979 32013 -973
rect 39107 -1013 39173 527
rect 39107 -1067 39113 -1013
rect 39167 -1067 39173 -1013
rect 39107 -1079 39173 -1067
rect 31867 -1131 32013 -1125
rect 21293 -1174 21462 -1168
rect 30252 -1174 30410 -1168
rect 14595 -1219 15439 -1216
rect 14593 -1282 15439 -1219
rect 14593 -2081 14659 -1282
rect 15373 -2081 15439 -1282
rect 14593 -2147 15439 -2081
<< via1 >>
rect 12978 4104 13030 4110
rect 12978 4040 13024 4104
rect 13024 4040 13030 4104
rect 12978 4034 13030 4040
rect 13574 4093 13626 4099
rect 13574 4053 13580 4093
rect 13580 4053 13620 4093
rect 13620 4053 13626 4093
rect 13574 4047 13626 4053
rect 14194 4093 14246 4099
rect 14194 4053 14200 4093
rect 14200 4053 14240 4093
rect 14240 4053 14246 4093
rect 14194 4047 14246 4053
rect 14834 4093 14886 4099
rect 14834 4053 14840 4093
rect 14840 4053 14880 4093
rect 14880 4053 14886 4093
rect 14834 4047 14886 4053
rect 15135 4047 15187 4099
rect 15454 4093 15506 4099
rect 15454 4053 15460 4093
rect 15460 4053 15500 4093
rect 15500 4053 15506 4093
rect 15454 4047 15506 4053
rect 16066 4104 16130 4110
rect 16066 4040 16124 4104
rect 16124 4040 16130 4104
rect 16066 4034 16130 4040
rect 16668 4098 16732 4104
rect 16668 4046 16674 4098
rect 16674 4046 16726 4098
rect 16726 4046 16732 4098
rect 16668 4040 16732 4046
rect 17048 4040 17112 4104
rect 17288 4098 17352 4104
rect 17288 4046 17294 4098
rect 17294 4046 17346 4098
rect 17346 4046 17352 4098
rect 17288 4040 17352 4046
rect 15786 3440 15792 3491
rect 15792 3440 15850 3491
rect 15850 3440 15856 3491
rect 15786 3434 15856 3440
rect 15136 2875 15188 2927
rect 14038 1744 14090 1750
rect 14038 1680 14084 1744
rect 14084 1680 14090 1744
rect 14038 1674 14090 1680
rect 14659 1744 14711 1750
rect 14659 1680 14665 1744
rect 14665 1680 14704 1744
rect 14704 1680 14711 1744
rect 14659 1674 14711 1680
rect 14954 1686 15006 1738
rect 15265 1744 15317 1750
rect 15265 1680 15272 1744
rect 15272 1680 15310 1744
rect 15310 1680 15317 1744
rect 15265 1674 15317 1680
rect 15886 1744 15938 1750
rect 15886 1680 15892 1744
rect 15892 1680 15938 1744
rect 15886 1674 15938 1680
rect 15606 1136 15674 1142
rect 15606 1086 15612 1136
rect 15612 1086 15668 1136
rect 15668 1086 15674 1136
rect 14954 494 15006 546
rect 17908 4098 17972 4104
rect 17908 4046 17914 4098
rect 17914 4046 17966 4098
rect 17966 4046 17972 4098
rect 17908 4040 17972 4046
rect 18528 4098 18592 4104
rect 18528 4046 18534 4098
rect 18534 4046 18586 4098
rect 18586 4046 18592 4098
rect 18528 4040 18592 4046
rect 19276 4104 19340 4110
rect 19276 4040 19334 4104
rect 19334 4040 19340 4104
rect 19276 4034 19340 4040
rect 19065 3432 19071 3485
rect 19071 3432 19131 3485
rect 19131 3432 19137 3485
rect 19065 3426 19137 3432
rect 17048 2228 17112 2292
rect 16512 1744 16564 1750
rect 16512 1680 16518 1744
rect 16518 1680 16561 1744
rect 16561 1680 16564 1744
rect 16512 1674 16564 1680
rect 17414 2876 17466 2928
rect 17409 2049 17472 2112
rect 34240 1752 34304 1758
rect 34240 1688 34298 1752
rect 34298 1688 34304 1752
rect 34240 1682 34304 1688
rect 17407 1487 17473 1553
rect 18486 1487 18552 1553
rect 25064 1336 25128 1342
rect 25064 1272 25070 1336
rect 25070 1272 25128 1336
rect 25064 1266 25128 1272
rect 26664 1336 26740 1342
rect 26664 1278 26670 1336
rect 26670 1278 26734 1336
rect 26734 1278 26740 1336
rect 20114 494 20166 546
rect 37118 527 37184 593
rect 39107 527 39173 593
rect 17048 -332 17112 -268
rect 18248 -332 18312 -268
rect 15618 -1073 15684 -1007
rect 17247 -1013 17313 -1007
rect 17247 -1067 17253 -1013
rect 17253 -1067 17307 -1013
rect 17307 -1067 17313 -1013
rect 17247 -1073 17313 -1067
rect 21305 -942 21462 -936
rect 21305 -1162 21456 -942
rect 21456 -1162 21462 -942
rect 21305 -1168 21462 -1162
rect 30264 -942 30410 -936
rect 22921 -979 23078 -973
rect 22921 -1124 22927 -979
rect 22927 -1124 23072 -979
rect 23072 -1124 23078 -979
rect 22921 -1130 23078 -1124
rect 30264 -1162 30404 -942
rect 30404 -1162 30410 -942
rect 30264 -1168 30410 -1162
rect 31867 -985 32013 -979
rect 31867 -1119 31873 -985
rect 31873 -1119 32007 -985
rect 32007 -1119 32013 -985
rect 31867 -1125 32013 -1119
<< metal2 >>
rect 12978 4110 13030 4116
rect 16066 4110 16130 4116
rect 19276 4110 19340 4116
rect 15135 4099 15187 4105
rect 13568 4098 13574 4099
rect 13030 4047 13574 4098
rect 13626 4098 13632 4099
rect 14188 4098 14194 4099
rect 13626 4047 14194 4098
rect 14246 4098 14252 4099
rect 14828 4098 14834 4099
rect 14246 4047 14834 4098
rect 14886 4098 14892 4099
rect 14886 4047 15135 4098
rect 15448 4098 15454 4099
rect 15187 4047 15454 4098
rect 15506 4047 15512 4099
rect 15135 4041 15187 4047
rect 12978 4028 13030 4034
rect 17048 4104 17112 4110
rect 16130 4040 16668 4104
rect 16732 4040 17048 4104
rect 17112 4040 17288 4104
rect 17352 4040 17908 4104
rect 17972 4040 18528 4104
rect 18592 4040 18598 4104
rect 17048 4034 17112 4040
rect 19340 4040 19726 4104
rect 16066 4028 16130 4034
rect 19276 4028 19340 4034
rect 15786 3493 15856 3502
rect 15780 3434 15786 3491
rect 15856 3434 15862 3491
rect 19065 3486 19137 3495
rect 15786 3424 15856 3433
rect 19059 3426 19065 3485
rect 19137 3426 19143 3485
rect 19065 3417 19137 3426
rect 20728 3372 20792 3381
rect 20728 3299 20792 3308
rect 15130 2924 15136 2927
rect 15120 2879 15136 2924
rect 15130 2875 15136 2879
rect 15188 2924 15194 2927
rect 17408 2924 17414 2928
rect 15188 2880 17414 2924
rect 15188 2875 15194 2880
rect 15460 2879 17414 2880
rect 17408 2876 17414 2879
rect 17466 2876 17472 2928
rect 17042 2228 17048 2292
rect 17112 2288 17852 2292
rect 17112 2232 17792 2288
rect 17848 2232 17857 2288
rect 17112 2228 17852 2232
rect 17654 2112 17710 2117
rect 17403 2049 17409 2112
rect 17472 2108 17714 2112
rect 17472 2052 17654 2108
rect 17710 2052 17714 2108
rect 17472 2049 17714 2052
rect 17654 2043 17710 2049
rect 34240 1758 34304 1764
rect 14038 1750 14090 1756
rect 14659 1750 14711 1756
rect 14090 1686 14659 1738
rect 14038 1668 14090 1674
rect 15265 1750 15317 1756
rect 14954 1738 15006 1744
rect 14711 1686 14954 1738
rect 15006 1686 15265 1738
rect 14954 1680 15006 1686
rect 14659 1668 14711 1674
rect 15886 1750 15938 1756
rect 15317 1686 15886 1738
rect 15265 1668 15317 1674
rect 16512 1750 16564 1756
rect 15938 1686 16512 1738
rect 15886 1668 15938 1674
rect 16564 1686 16586 1738
rect 34304 1688 34708 1752
rect 34240 1676 34304 1682
rect 16512 1668 16564 1674
rect 17407 1553 17473 1559
rect 18486 1553 18552 1559
rect 17473 1487 18486 1553
rect 17407 1481 17473 1487
rect 18486 1481 18552 1487
rect 25064 1342 25128 1348
rect 26664 1342 26740 1351
rect 25055 1266 25064 1342
rect 25128 1266 25137 1342
rect 26658 1278 26664 1342
rect 26740 1278 26746 1342
rect 26664 1269 26740 1278
rect 25064 1260 25128 1266
rect 15606 1144 15674 1153
rect 15600 1086 15606 1142
rect 15674 1086 15680 1142
rect 15606 1075 15674 1084
rect 14954 546 15006 552
rect 20114 546 20166 552
rect 15006 494 20114 546
rect 20166 494 20186 546
rect 37107 527 37118 593
rect 37184 527 39107 593
rect 39173 527 39179 593
rect 14954 488 15006 494
rect 20114 488 20166 494
rect 17048 -268 17112 -262
rect 18248 -268 18312 -262
rect 17112 -332 18248 -268
rect 17048 -338 17112 -332
rect 18248 -338 18312 -332
rect 21305 -936 21462 -930
rect 15618 -1007 15684 -1001
rect 17247 -1007 17313 -1001
rect 15684 -1073 17247 -1007
rect 15618 -1079 15684 -1073
rect 17247 -1079 17313 -1073
rect 30264 -936 30410 -930
rect 21462 -1130 22921 -973
rect 23078 -1130 23084 -973
rect 21305 -1174 21462 -1168
rect 30410 -1125 31867 -979
rect 32013 -1125 32019 -979
rect 30264 -1174 30410 -1168
<< via2 >>
rect 15786 3491 15856 3493
rect 15786 3434 15856 3491
rect 19065 3485 19137 3486
rect 15786 3433 15856 3434
rect 19065 3426 19137 3485
rect 20728 3308 20792 3372
rect 17792 2232 17848 2288
rect 17654 2052 17710 2108
rect 25064 1266 25128 1342
rect 26664 1278 26740 1342
rect 15606 1142 15674 1144
rect 15606 1086 15674 1142
rect 15606 1084 15674 1086
<< metal3 >>
rect 15781 3493 15861 3498
rect 15781 3433 15786 3493
rect 15856 3433 15861 3493
rect 15781 3428 15861 3433
rect 19060 3486 19142 3491
rect 15791 3280 15851 3428
rect 19060 3426 19065 3486
rect 19137 3426 19142 3486
rect 19060 3421 19142 3426
rect 15790 3230 15851 3280
rect 15790 2798 15850 3230
rect 15608 2792 15672 2798
rect 15608 2722 15672 2728
rect 15788 2792 15852 2798
rect 19071 2792 19131 3421
rect 20723 3372 20797 3377
rect 20723 3308 20728 3372
rect 20792 3308 20797 3372
rect 20723 3303 20797 3308
rect 20728 2792 20792 3303
rect 19063 2728 19069 2792
rect 19133 2728 19139 2792
rect 20722 2728 20728 2792
rect 20792 2728 20798 2792
rect 15788 2722 15852 2728
rect 15610 1149 15670 2722
rect 17787 2288 17853 2293
rect 17787 2232 17792 2288
rect 17848 2232 17853 2288
rect 17787 2227 17853 2232
rect 17649 2108 17715 2113
rect 17788 2112 17852 2227
rect 17649 2052 17654 2108
rect 17710 2052 17715 2108
rect 17649 2047 17715 2052
rect 17782 2048 17788 2112
rect 17852 2048 17858 2112
rect 26664 2048 26670 2112
rect 26734 2048 26740 2112
rect 17650 1959 17713 2047
rect 17649 1953 17713 1959
rect 17649 1883 17713 1889
rect 25058 1888 25064 1952
rect 25128 1888 25134 1952
rect 25064 1347 25128 1888
rect 26670 1347 26734 2048
rect 25059 1342 25133 1347
rect 25059 1266 25064 1342
rect 25128 1266 25133 1342
rect 26659 1342 26745 1347
rect 26659 1278 26664 1342
rect 26740 1278 26745 1342
rect 26659 1273 26745 1278
rect 25059 1261 25133 1266
rect 15601 1144 15679 1149
rect 15601 1084 15606 1144
rect 15674 1084 15679 1144
rect 15601 1079 15679 1084
<< via3 >>
rect 15608 2728 15672 2792
rect 15788 2728 15852 2792
rect 19069 2728 19133 2792
rect 20728 2728 20792 2792
rect 17788 2048 17852 2112
rect 26670 2048 26734 2112
rect 17649 1889 17713 1953
rect 25064 1888 25128 1952
<< metal4 >>
rect 15607 2792 15673 2793
rect 15787 2792 15853 2793
rect 19068 2792 19134 2793
rect 20727 2792 20793 2793
rect 15460 2728 15608 2792
rect 15672 2728 15788 2792
rect 15852 2728 19069 2792
rect 19133 2728 20728 2792
rect 20792 2728 20793 2792
rect 15607 2727 15673 2728
rect 15787 2727 15853 2728
rect 19068 2727 19134 2728
rect 20727 2727 20793 2728
rect 17787 2112 17853 2113
rect 26669 2112 26735 2113
rect 17787 2048 17788 2112
rect 17852 2048 26670 2112
rect 26734 2048 26735 2112
rect 17787 2047 17853 2048
rect 26669 2047 26735 2048
rect 17648 1953 17714 1954
rect 17648 1889 17649 1953
rect 17713 1952 17714 1953
rect 25063 1952 25129 1953
rect 17713 1889 25064 1952
rect 17648 1888 17714 1889
rect 24248 1888 25064 1889
rect 25128 1888 25129 1952
rect 25063 1887 25129 1888
use CM_OTA_NCH  CM_OTA_NCH_0
timestamp 1711300264
transform -1 0 27500 0 1 900
box -7620 -1100 8200 5936
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 13984 -1 0 4872
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_1
timestamp 1695852000
transform 0 1 12744 -1 0 4872
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_2
timestamp 1695852000
transform 0 1 13364 -1 0 4872
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_4
timestamp 1695852000
transform 0 1 18324 -1 0 4872
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_13
timestamp 1695852000
transform 0 1 15684 -1 0 2512
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_19
timestamp 1695852000
transform 0 1 15064 -1 0 2512
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_20
timestamp 1695852000
transform 0 1 15224 -1 0 4872
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_35
timestamp 1695852000
transform 0 1 14424 -1 0 2512
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_37
timestamp 1695852000
transform 0 1 13804 -1 0 2512
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_39
timestamp 1695852000
transform 0 1 14604 -1 0 4872
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_41
timestamp 1695852000
transform 0 1 16310 -1 0 2512
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_59
timestamp 1695852000
transform 0 1 17084 -1 0 4872
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_60
timestamp 1695852000
transform 0 1 17704 -1 0 4872
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_61
timestamp 1695852000
transform 0 1 15844 -1 0 4872
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_62
timestamp 1695852000
transform 0 1 16464 -1 0 4872
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_63
timestamp 1695852000
transform 0 1 19060 -1 0 4872
box -184 -124 1912 613
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 1 1288 0 1 1288
timestamp 1704988097
transform 1 0 35200 0 1 820
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1704988097
transform 1 0 17856 0 1 860
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_2
array 0 1 1288 0 1 1288
timestamp 1704988097
transform 1 0 13700 0 1 -3000
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_3
timestamp 1704988097
transform 1 0 37840 0 1 820
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_4
timestamp 1704988097
transform 1 0 12340 0 1 -1720
box 0 0 1340 1340
use SUNTR_RPPO2  SUNTR_RPPO2_0 ~/aicex/ip/cnr_gr03_sky130nm/design/SUN_TR_SKY130NM
timestamp 1710432512
transform 1 0 16500 0 1 -4600
box 0 0 2672 4236
use SUNTR_RPPO2  SUNTR_RPPO2_1
timestamp 1710432512
transform -1 0 22072 0 1 -4600
box 0 0 2672 4236
use SUNTR_RPPO16  SUNTR_RPPO16_0 ~/aicex/ip/cnr_gr03_sky130nm/design/SUN_TR_SKY130NM
timestamp 1710432512
transform -1 0 39920 0 1 -4600
box 0 0 8720 4236
use SUNTR_RPPO16  SUNTR_RPPO16_1
timestamp 1710432512
transform -1 0 31020 0 1 -4600
box 0 0 8720 4236
<< labels >>
flabel locali 16326 -200 19500 0 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel locali 14100 160 19230 360 0 FreeSans 800 0 0 0 VSS
port 4 nsew
flabel metal2 19340 4040 19726 4104 0 FreeSans 1600 0 0 0 I_OUT1
port 9 nsew
flabel metal2 15006 494 20114 546 0 FreeSans 800 0 0 0 VREF
port 10 nsew
flabel metal2 34304 1688 34708 1752 0 FreeSans 800 0 0 0 IBIAS
port 7 nsew
flabel space 17409 1227 17471 2876 0 FreeSans 800 0 0 0 VD1
flabel metal1 17048 -268 17112 4030 0 FreeSans 800 0 0 0 VR1
<< end >>

