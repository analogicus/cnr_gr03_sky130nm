*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/MILESTONE2_lpe.spi
#else
.include ../../../work/xsch/MILESTONE2.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0 dc 0
VDD  VDD_1V8 VSS dc 1.8
VRST RST VSS PULSE(0 1.8 0.0 2NS 2NS 75NS 275NS)
*VRST RST VSS dc 0
IIN VSS I_IN dc 60u
VREF VREF_I VSS dc 1.2

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT RST OUT I_IN VREF_I VDD_1V8 VSS MILESTONE2

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save v(OUT) v(VDD) v(VSS) v(RST) v(VREF_I) v(I_IN) 
*.save all
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquitex

optran 0 0 0 10n 10u 0
tran 1n 1u 0.3u
write {cicname}_tran.raw


*dc IIN 50u 75u 100n
write
quit

.endc

.end
