magic
tech sky130B
magscale 1 2
timestamp 1712935398
<< viali >>
rect 6561 9605 6595 9639
rect 6377 9401 6411 9435
rect 7389 9061 7423 9095
rect 8677 9061 8711 9095
rect 6009 8993 6043 9027
rect 7757 8993 7791 9027
rect 8033 8993 8067 9027
rect 1961 8925 1995 8959
rect 4353 8925 4387 8959
rect 4537 8925 4571 8959
rect 7665 8925 7699 8959
rect 8493 8925 8527 8959
rect 2228 8857 2262 8891
rect 4804 8857 4838 8891
rect 6254 8857 6288 8891
rect 3341 8789 3375 8823
rect 3801 8789 3835 8823
rect 5917 8789 5951 8823
rect 2973 8585 3007 8619
rect 5733 8585 5767 8619
rect 6622 8517 6656 8551
rect 1676 8449 1710 8483
rect 2881 8449 2915 8483
rect 3065 8449 3099 8483
rect 3157 8449 3191 8483
rect 5917 8449 5951 8483
rect 6377 8449 6411 8483
rect 1409 8381 1443 8415
rect 5549 8381 5583 8415
rect 2789 8245 2823 8279
rect 4629 8245 4663 8279
rect 4997 8245 5031 8279
rect 7757 8245 7791 8279
rect 2053 8041 2087 8075
rect 5549 8041 5583 8075
rect 1593 7973 1627 8007
rect 5181 7973 5215 8007
rect 3617 7905 3651 7939
rect 1409 7837 1443 7871
rect 2237 7837 2271 7871
rect 2513 7837 2547 7871
rect 3249 7837 3283 7871
rect 3341 7837 3375 7871
rect 3433 7837 3467 7871
rect 3808 7837 3842 7871
rect 5549 7837 5583 7871
rect 5641 7837 5675 7871
rect 5825 7837 5859 7871
rect 8493 7837 8527 7871
rect 4046 7769 4080 7803
rect 2421 7701 2455 7735
rect 2605 7701 2639 7735
rect 3617 7701 3651 7735
rect 5365 7701 5399 7735
rect 8677 7701 8711 7735
rect 2329 7497 2363 7531
rect 2697 7497 2731 7531
rect 3525 7497 3559 7531
rect 7849 7497 7883 7531
rect 8125 7497 8159 7531
rect 2605 7361 2639 7395
rect 2881 7361 2915 7395
rect 2973 7361 3007 7395
rect 3157 7361 3191 7395
rect 4077 7361 4111 7395
rect 4353 7361 4387 7395
rect 4629 7361 4663 7395
rect 5457 7361 5491 7395
rect 5733 7361 5767 7395
rect 6009 7361 6043 7395
rect 6377 7361 6411 7395
rect 6633 7361 6667 7395
rect 8033 7361 8067 7395
rect 8217 7361 8251 7395
rect 2329 7293 2363 7327
rect 3801 7293 3835 7327
rect 4445 7293 4479 7327
rect 4537 7293 4571 7327
rect 5825 7293 5859 7327
rect 2513 7225 2547 7259
rect 3065 7225 3099 7259
rect 8401 7225 8435 7259
rect 3985 7157 4019 7191
rect 4169 7157 4203 7191
rect 4813 7157 4847 7191
rect 5549 7157 5583 7191
rect 5733 7157 5767 7191
rect 7757 7157 7791 7191
rect 4077 6953 4111 6987
rect 7481 6885 7515 6919
rect 7849 6817 7883 6851
rect 8125 6817 8159 6851
rect 8401 6817 8435 6851
rect 2881 6749 2915 6783
rect 3433 6749 3467 6783
rect 3617 6749 3651 6783
rect 3801 6749 3835 6783
rect 4261 6749 4295 6783
rect 4353 6749 4387 6783
rect 4537 6749 4571 6783
rect 4629 6749 4663 6783
rect 5549 6749 5583 6783
rect 7205 6749 7239 6783
rect 7757 6749 7791 6783
rect 2614 6681 2648 6715
rect 3525 6681 3559 6715
rect 5816 6681 5850 6715
rect 7481 6681 7515 6715
rect 8677 6681 8711 6715
rect 1501 6613 1535 6647
rect 3893 6613 3927 6647
rect 6929 6613 6963 6647
rect 7297 6613 7331 6647
rect 6009 6409 6043 6443
rect 8769 6409 8803 6443
rect 8217 6341 8251 6375
rect 8417 6341 8451 6375
rect 1777 6273 1811 6307
rect 2973 6273 3007 6307
rect 3433 6273 3467 6307
rect 3985 6273 4019 6307
rect 4344 6273 4378 6307
rect 6193 6273 6227 6307
rect 7573 6273 7607 6307
rect 8677 6273 8711 6307
rect 8861 6273 8895 6307
rect 4077 6205 4111 6239
rect 7665 6205 7699 6239
rect 3157 6137 3191 6171
rect 5457 6137 5491 6171
rect 8585 6137 8619 6171
rect 2421 6069 2455 6103
rect 2697 6069 2731 6103
rect 3065 6069 3099 6103
rect 3249 6069 3283 6103
rect 3801 6069 3835 6103
rect 7941 6069 7975 6103
rect 8401 6069 8435 6103
rect 1501 5865 1535 5899
rect 2421 5865 2455 5899
rect 5089 5865 5123 5899
rect 8677 5865 8711 5899
rect 2789 5797 2823 5831
rect 2513 5729 2547 5763
rect 1777 5661 1811 5695
rect 2145 5661 2179 5695
rect 2237 5661 2271 5695
rect 2329 5661 2363 5695
rect 2605 5661 2639 5695
rect 2881 5661 2915 5695
rect 3801 5661 3835 5695
rect 6193 5661 6227 5695
rect 7665 5661 7699 5695
rect 7849 5661 7883 5695
rect 8493 5661 8527 5695
rect 2053 5593 2087 5627
rect 2881 5525 2915 5559
rect 5641 5525 5675 5559
rect 7757 5525 7791 5559
rect 3709 5321 3743 5355
rect 4077 5321 4111 5355
rect 2145 5185 2179 5219
rect 2237 5185 2271 5219
rect 2421 5185 2455 5219
rect 2513 5185 2547 5219
rect 3341 5185 3375 5219
rect 3525 5185 3559 5219
rect 3985 5185 4019 5219
rect 4169 5185 4203 5219
rect 4712 5185 4746 5219
rect 6633 5185 6667 5219
rect 8033 5185 8067 5219
rect 8585 5185 8619 5219
rect 2605 5117 2639 5151
rect 3157 5117 3191 5151
rect 4445 5117 4479 5151
rect 6377 5117 6411 5151
rect 7941 5117 7975 5151
rect 1961 4981 1995 5015
rect 5825 4981 5859 5015
rect 7757 4981 7791 5015
rect 8309 4981 8343 5015
rect 8769 4981 8803 5015
rect 2789 4777 2823 4811
rect 3249 4777 3283 4811
rect 3985 4777 4019 4811
rect 4261 4777 4295 4811
rect 4537 4777 4571 4811
rect 5273 4777 5307 4811
rect 7573 4777 7607 4811
rect 3801 4709 3835 4743
rect 5089 4709 5123 4743
rect 7021 4709 7055 4743
rect 7389 4641 7423 4675
rect 1409 4573 1443 4607
rect 1676 4573 1710 4607
rect 3065 4573 3099 4607
rect 3341 4573 3375 4607
rect 3985 4573 4019 4607
rect 4169 4573 4203 4607
rect 4445 4573 4479 4607
rect 4537 4573 4571 4607
rect 4721 4573 4755 4607
rect 4813 4573 4847 4607
rect 5089 4573 5123 4607
rect 5181 4573 5215 4607
rect 5365 4573 5399 4607
rect 5641 4573 5675 4607
rect 7297 4573 7331 4607
rect 7757 4573 7791 4607
rect 8033 4573 8067 4607
rect 8217 4573 8251 4607
rect 8493 4573 8527 4607
rect 5886 4505 5920 4539
rect 2881 4437 2915 4471
rect 4905 4437 4939 4471
rect 8677 4437 8711 4471
rect 2789 4097 2823 4131
rect 5181 4097 5215 4131
rect 7481 4097 7515 4131
rect 7665 4097 7699 4131
rect 7757 4097 7791 4131
rect 7849 4097 7883 4131
rect 2513 4029 2547 4063
rect 4905 4029 4939 4063
rect 8125 4029 8159 4063
rect 2237 3893 2271 3927
rect 2697 3893 2731 3927
rect 4997 3893 5031 3927
rect 5089 3893 5123 3927
rect 4629 3689 4663 3723
rect 5181 3689 5215 3723
rect 4813 3621 4847 3655
rect 8677 3621 8711 3655
rect 4353 3553 4387 3587
rect 4537 3553 4571 3587
rect 5733 3553 5767 3587
rect 1961 3485 1995 3519
rect 4077 3485 4111 3519
rect 4261 3485 4295 3519
rect 4445 3485 4479 3519
rect 5917 3485 5951 3519
rect 7849 3485 7883 3519
rect 8033 3485 8067 3519
rect 8493 3485 8527 3519
rect 6162 3417 6196 3451
rect 1777 3349 1811 3383
rect 3893 3349 3927 3383
rect 7297 3349 7331 3383
rect 7941 3349 7975 3383
rect 2789 3145 2823 3179
rect 6101 3145 6135 3179
rect 7757 3145 7791 3179
rect 4629 3077 4663 3111
rect 6622 3077 6656 3111
rect 8217 3077 8251 3111
rect 8493 3077 8527 3111
rect 1409 3009 1443 3043
rect 1676 3009 1710 3043
rect 4988 3009 5022 3043
rect 6377 3009 6411 3043
rect 8033 3009 8067 3043
rect 8309 3009 8343 3043
rect 4721 2941 4755 2975
rect 7849 2941 7883 2975
rect 3341 2873 3375 2907
rect 8677 2805 8711 2839
rect 3617 2601 3651 2635
rect 4353 2601 4387 2635
rect 4629 2601 4663 2635
rect 8033 2601 8067 2635
rect 8677 2601 8711 2635
rect 3893 2533 3927 2567
rect 2237 2465 2271 2499
rect 1961 2397 1995 2431
rect 4169 2397 4203 2431
rect 4445 2397 4479 2431
rect 4905 2397 4939 2431
rect 7665 2397 7699 2431
rect 7941 2397 7975 2431
rect 2482 2329 2516 2363
rect 4629 2329 4663 2363
rect 4813 2329 4847 2363
rect 8401 2329 8435 2363
rect 2145 2261 2179 2295
rect 7849 2261 7883 2295
<< metal1 >>
rect 1104 9818 9200 9840
rect 1104 9766 2622 9818
rect 2674 9766 2686 9818
rect 2738 9766 2750 9818
rect 2802 9766 2814 9818
rect 2866 9766 2878 9818
rect 2930 9766 4646 9818
rect 4698 9766 4710 9818
rect 4762 9766 4774 9818
rect 4826 9766 4838 9818
rect 4890 9766 4902 9818
rect 4954 9766 6670 9818
rect 6722 9766 6734 9818
rect 6786 9766 6798 9818
rect 6850 9766 6862 9818
rect 6914 9766 6926 9818
rect 6978 9766 8694 9818
rect 8746 9766 8758 9818
rect 8810 9766 8822 9818
rect 8874 9766 8886 9818
rect 8938 9766 8950 9818
rect 9002 9766 9200 9818
rect 1104 9744 9200 9766
rect 5810 9596 5816 9648
rect 5868 9636 5874 9648
rect 6549 9639 6607 9645
rect 6549 9636 6561 9639
rect 5868 9608 6561 9636
rect 5868 9596 5874 9608
rect 6549 9605 6561 9608
rect 6595 9605 6607 9639
rect 6549 9599 6607 9605
rect 6362 9392 6368 9444
rect 6420 9392 6426 9444
rect 1104 9274 9200 9296
rect 1104 9222 1962 9274
rect 2014 9222 2026 9274
rect 2078 9222 2090 9274
rect 2142 9222 2154 9274
rect 2206 9222 2218 9274
rect 2270 9222 3986 9274
rect 4038 9222 4050 9274
rect 4102 9222 4114 9274
rect 4166 9222 4178 9274
rect 4230 9222 4242 9274
rect 4294 9222 6010 9274
rect 6062 9222 6074 9274
rect 6126 9222 6138 9274
rect 6190 9222 6202 9274
rect 6254 9222 6266 9274
rect 6318 9222 8034 9274
rect 8086 9222 8098 9274
rect 8150 9222 8162 9274
rect 8214 9222 8226 9274
rect 8278 9222 8290 9274
rect 8342 9222 9200 9274
rect 1104 9200 9200 9222
rect 6362 9160 6368 9172
rect 6012 9132 6368 9160
rect 6012 9033 6040 9132
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 7377 9095 7435 9101
rect 7377 9061 7389 9095
rect 7423 9061 7435 9095
rect 7377 9055 7435 9061
rect 5997 9027 6055 9033
rect 5997 8993 6009 9027
rect 6043 8993 6055 9027
rect 5997 8987 6055 8993
rect 1486 8916 1492 8968
rect 1544 8956 1550 8968
rect 1949 8959 2007 8965
rect 1949 8956 1961 8959
rect 1544 8928 1961 8956
rect 1544 8916 1550 8928
rect 1949 8925 1961 8928
rect 1995 8956 2007 8959
rect 1995 8928 3372 8956
rect 1995 8925 2007 8928
rect 1949 8919 2007 8925
rect 2216 8891 2274 8897
rect 2216 8857 2228 8891
rect 2262 8888 2274 8891
rect 2958 8888 2964 8900
rect 2262 8860 2964 8888
rect 2262 8857 2274 8860
rect 2216 8851 2274 8857
rect 2958 8848 2964 8860
rect 3016 8848 3022 8900
rect 3344 8888 3372 8928
rect 4338 8916 4344 8968
rect 4396 8916 4402 8968
rect 4522 8916 4528 8968
rect 4580 8916 4586 8968
rect 7392 8956 7420 9055
rect 8662 9052 8668 9104
rect 8720 9052 8726 9104
rect 7742 8984 7748 9036
rect 7800 8984 7806 9036
rect 8021 9027 8079 9033
rect 8021 8993 8033 9027
rect 8067 9024 8079 9027
rect 8067 8996 8524 9024
rect 8067 8993 8079 8996
rect 8021 8987 8079 8993
rect 8496 8965 8524 8996
rect 7653 8959 7711 8965
rect 7653 8956 7665 8959
rect 7392 8928 7665 8956
rect 7653 8925 7665 8928
rect 7699 8925 7711 8959
rect 7653 8919 7711 8925
rect 8481 8959 8539 8965
rect 8481 8925 8493 8959
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 4540 8888 4568 8916
rect 3344 8860 4568 8888
rect 4792 8891 4850 8897
rect 4792 8857 4804 8891
rect 4838 8888 4850 8891
rect 5718 8888 5724 8900
rect 4838 8860 5724 8888
rect 4838 8857 4850 8860
rect 4792 8851 4850 8857
rect 5718 8848 5724 8860
rect 5776 8848 5782 8900
rect 5810 8848 5816 8900
rect 5868 8888 5874 8900
rect 6242 8891 6300 8897
rect 6242 8888 6254 8891
rect 5868 8860 6254 8888
rect 5868 8848 5874 8860
rect 6242 8857 6254 8860
rect 6288 8857 6300 8891
rect 6242 8851 6300 8857
rect 3050 8780 3056 8832
rect 3108 8820 3114 8832
rect 3329 8823 3387 8829
rect 3329 8820 3341 8823
rect 3108 8792 3341 8820
rect 3108 8780 3114 8792
rect 3329 8789 3341 8792
rect 3375 8789 3387 8823
rect 3329 8783 3387 8789
rect 3418 8780 3424 8832
rect 3476 8820 3482 8832
rect 3789 8823 3847 8829
rect 3789 8820 3801 8823
rect 3476 8792 3801 8820
rect 3476 8780 3482 8792
rect 3789 8789 3801 8792
rect 3835 8789 3847 8823
rect 3789 8783 3847 8789
rect 5626 8780 5632 8832
rect 5684 8820 5690 8832
rect 5905 8823 5963 8829
rect 5905 8820 5917 8823
rect 5684 8792 5917 8820
rect 5684 8780 5690 8792
rect 5905 8789 5917 8792
rect 5951 8789 5963 8823
rect 5905 8783 5963 8789
rect 1104 8730 9200 8752
rect 1104 8678 2622 8730
rect 2674 8678 2686 8730
rect 2738 8678 2750 8730
rect 2802 8678 2814 8730
rect 2866 8678 2878 8730
rect 2930 8678 4646 8730
rect 4698 8678 4710 8730
rect 4762 8678 4774 8730
rect 4826 8678 4838 8730
rect 4890 8678 4902 8730
rect 4954 8678 6670 8730
rect 6722 8678 6734 8730
rect 6786 8678 6798 8730
rect 6850 8678 6862 8730
rect 6914 8678 6926 8730
rect 6978 8678 8694 8730
rect 8746 8678 8758 8730
rect 8810 8678 8822 8730
rect 8874 8678 8886 8730
rect 8938 8678 8950 8730
rect 9002 8678 9200 8730
rect 1104 8656 9200 8678
rect 2958 8576 2964 8628
rect 3016 8576 3022 8628
rect 3418 8576 3424 8628
rect 3476 8576 3482 8628
rect 5718 8576 5724 8628
rect 5776 8576 5782 8628
rect 3436 8548 3464 8576
rect 6610 8551 6668 8557
rect 6610 8548 6622 8551
rect 3068 8520 3464 8548
rect 5644 8520 6622 8548
rect 1486 8480 1492 8492
rect 1412 8452 1492 8480
rect 1412 8421 1440 8452
rect 1486 8440 1492 8452
rect 1544 8440 1550 8492
rect 1670 8489 1676 8492
rect 1664 8443 1676 8489
rect 1670 8440 1676 8443
rect 1728 8440 1734 8492
rect 2498 8440 2504 8492
rect 2556 8480 2562 8492
rect 3068 8489 3096 8520
rect 5644 8492 5672 8520
rect 6610 8517 6622 8520
rect 6656 8517 6668 8551
rect 6610 8511 6668 8517
rect 2869 8483 2927 8489
rect 2869 8480 2881 8483
rect 2556 8452 2881 8480
rect 2556 8440 2562 8452
rect 2869 8449 2881 8452
rect 2915 8449 2927 8483
rect 2869 8443 2927 8449
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8480 3203 8483
rect 5074 8480 5080 8492
rect 3191 8452 5080 8480
rect 3191 8449 3203 8452
rect 3145 8443 3203 8449
rect 5074 8440 5080 8452
rect 5132 8440 5138 8492
rect 5626 8440 5632 8492
rect 5684 8440 5690 8492
rect 5718 8440 5724 8492
rect 5776 8480 5782 8492
rect 5905 8483 5963 8489
rect 5905 8480 5917 8483
rect 5776 8452 5917 8480
rect 5776 8440 5782 8452
rect 5905 8449 5917 8452
rect 5951 8449 5963 8483
rect 5905 8443 5963 8449
rect 6362 8440 6368 8492
rect 6420 8440 6426 8492
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8381 1455 8415
rect 1397 8375 1455 8381
rect 5534 8372 5540 8424
rect 5592 8372 5598 8424
rect 2777 8279 2835 8285
rect 2777 8245 2789 8279
rect 2823 8276 2835 8279
rect 3234 8276 3240 8288
rect 2823 8248 3240 8276
rect 2823 8245 2835 8248
rect 2777 8239 2835 8245
rect 3234 8236 3240 8248
rect 3292 8236 3298 8288
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 4522 8276 4528 8288
rect 3476 8248 4528 8276
rect 3476 8236 3482 8248
rect 4522 8236 4528 8248
rect 4580 8236 4586 8288
rect 4614 8236 4620 8288
rect 4672 8236 4678 8288
rect 4982 8236 4988 8288
rect 5040 8236 5046 8288
rect 7745 8279 7803 8285
rect 7745 8245 7757 8279
rect 7791 8276 7803 8279
rect 7926 8276 7932 8288
rect 7791 8248 7932 8276
rect 7791 8245 7803 8248
rect 7745 8239 7803 8245
rect 7926 8236 7932 8248
rect 7984 8236 7990 8288
rect 1104 8186 9200 8208
rect 1104 8134 1962 8186
rect 2014 8134 2026 8186
rect 2078 8134 2090 8186
rect 2142 8134 2154 8186
rect 2206 8134 2218 8186
rect 2270 8134 3986 8186
rect 4038 8134 4050 8186
rect 4102 8134 4114 8186
rect 4166 8134 4178 8186
rect 4230 8134 4242 8186
rect 4294 8134 6010 8186
rect 6062 8134 6074 8186
rect 6126 8134 6138 8186
rect 6190 8134 6202 8186
rect 6254 8134 6266 8186
rect 6318 8134 8034 8186
rect 8086 8134 8098 8186
rect 8150 8134 8162 8186
rect 8214 8134 8226 8186
rect 8278 8134 8290 8186
rect 8342 8134 9200 8186
rect 1104 8112 9200 8134
rect 1670 8032 1676 8084
rect 1728 8072 1734 8084
rect 2041 8075 2099 8081
rect 2041 8072 2053 8075
rect 1728 8044 2053 8072
rect 1728 8032 1734 8044
rect 2041 8041 2053 8044
rect 2087 8041 2099 8075
rect 4982 8072 4988 8084
rect 2041 8035 2099 8041
rect 3620 8044 4988 8072
rect 1581 8007 1639 8013
rect 1581 7973 1593 8007
rect 1627 8004 1639 8007
rect 3510 8004 3516 8016
rect 1627 7976 3516 8004
rect 1627 7973 1639 7976
rect 1581 7967 1639 7973
rect 3510 7964 3516 7976
rect 3568 7964 3574 8016
rect 3620 7945 3648 8044
rect 4982 8032 4988 8044
rect 5040 8032 5046 8084
rect 5534 8032 5540 8084
rect 5592 8032 5598 8084
rect 5169 8007 5227 8013
rect 5169 7973 5181 8007
rect 5215 8004 5227 8007
rect 5215 7976 5856 8004
rect 5215 7973 5227 7976
rect 5169 7967 5227 7973
rect 3605 7939 3663 7945
rect 2746 7908 3464 7936
rect 1394 7828 1400 7880
rect 1452 7828 1458 7880
rect 2222 7828 2228 7880
rect 2280 7828 2286 7880
rect 2501 7871 2559 7877
rect 2501 7837 2513 7871
rect 2547 7868 2559 7871
rect 2746 7868 2774 7908
rect 3436 7880 3464 7908
rect 3605 7905 3617 7939
rect 3651 7905 3663 7939
rect 3605 7899 3663 7905
rect 5828 7880 5856 7976
rect 2547 7840 2774 7868
rect 2547 7837 2559 7840
rect 2501 7831 2559 7837
rect 3234 7828 3240 7880
rect 3292 7868 3298 7880
rect 3329 7871 3387 7877
rect 3329 7868 3341 7871
rect 3292 7840 3341 7868
rect 3292 7828 3298 7840
rect 3329 7837 3341 7840
rect 3375 7837 3387 7871
rect 3329 7831 3387 7837
rect 3344 7800 3372 7831
rect 3418 7828 3424 7880
rect 3476 7828 3482 7880
rect 3510 7828 3516 7880
rect 3568 7828 3574 7880
rect 3796 7871 3854 7877
rect 3796 7837 3808 7871
rect 3842 7868 3854 7871
rect 4614 7868 4620 7880
rect 3842 7840 4620 7868
rect 3842 7837 3854 7840
rect 3796 7831 3854 7837
rect 3528 7800 3556 7828
rect 4172 7812 4200 7840
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 5537 7871 5595 7877
rect 5537 7837 5549 7871
rect 5583 7837 5595 7871
rect 5537 7831 5595 7837
rect 3344 7772 3556 7800
rect 3694 7760 3700 7812
rect 3752 7800 3758 7812
rect 4034 7803 4092 7809
rect 4034 7800 4046 7803
rect 3752 7772 4046 7800
rect 3752 7760 3758 7772
rect 4034 7769 4046 7772
rect 4080 7769 4092 7803
rect 4034 7763 4092 7769
rect 4154 7760 4160 7812
rect 4212 7760 4218 7812
rect 4338 7760 4344 7812
rect 4396 7760 4402 7812
rect 4430 7760 4436 7812
rect 4488 7800 4494 7812
rect 5552 7800 5580 7831
rect 5626 7828 5632 7880
rect 5684 7828 5690 7880
rect 5810 7828 5816 7880
rect 5868 7828 5874 7880
rect 5902 7828 5908 7880
rect 5960 7828 5966 7880
rect 8478 7828 8484 7880
rect 8536 7828 8542 7880
rect 5920 7800 5948 7828
rect 4488 7772 5948 7800
rect 4488 7760 4494 7772
rect 2409 7735 2467 7741
rect 2409 7701 2421 7735
rect 2455 7732 2467 7735
rect 2593 7735 2651 7741
rect 2593 7732 2605 7735
rect 2455 7704 2605 7732
rect 2455 7701 2467 7704
rect 2409 7695 2467 7701
rect 2593 7701 2605 7704
rect 2639 7701 2651 7735
rect 2593 7695 2651 7701
rect 3605 7735 3663 7741
rect 3605 7701 3617 7735
rect 3651 7732 3663 7735
rect 4356 7732 4384 7760
rect 3651 7704 4384 7732
rect 3651 7701 3663 7704
rect 3605 7695 3663 7701
rect 5350 7692 5356 7744
rect 5408 7692 5414 7744
rect 8665 7735 8723 7741
rect 8665 7701 8677 7735
rect 8711 7732 8723 7735
rect 9122 7732 9128 7744
rect 8711 7704 9128 7732
rect 8711 7701 8723 7704
rect 8665 7695 8723 7701
rect 9122 7692 9128 7704
rect 9180 7692 9186 7744
rect 1104 7642 9200 7664
rect 1104 7590 2622 7642
rect 2674 7590 2686 7642
rect 2738 7590 2750 7642
rect 2802 7590 2814 7642
rect 2866 7590 2878 7642
rect 2930 7590 4646 7642
rect 4698 7590 4710 7642
rect 4762 7590 4774 7642
rect 4826 7590 4838 7642
rect 4890 7590 4902 7642
rect 4954 7590 6670 7642
rect 6722 7590 6734 7642
rect 6786 7590 6798 7642
rect 6850 7590 6862 7642
rect 6914 7590 6926 7642
rect 6978 7590 8694 7642
rect 8746 7590 8758 7642
rect 8810 7590 8822 7642
rect 8874 7590 8886 7642
rect 8938 7590 8950 7642
rect 9002 7590 9200 7642
rect 1104 7568 9200 7590
rect 2222 7488 2228 7540
rect 2280 7528 2286 7540
rect 2317 7531 2375 7537
rect 2317 7528 2329 7531
rect 2280 7500 2329 7528
rect 2280 7488 2286 7500
rect 2317 7497 2329 7500
rect 2363 7497 2375 7531
rect 2317 7491 2375 7497
rect 2498 7488 2504 7540
rect 2556 7528 2562 7540
rect 2685 7531 2743 7537
rect 2685 7528 2697 7531
rect 2556 7500 2697 7528
rect 2556 7488 2562 7500
rect 2685 7497 2697 7500
rect 2731 7497 2743 7531
rect 3234 7528 3240 7540
rect 2685 7491 2743 7497
rect 2884 7500 3240 7528
rect 2884 7401 2912 7500
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 3513 7531 3571 7537
rect 3513 7497 3525 7531
rect 3559 7528 3571 7531
rect 5718 7528 5724 7540
rect 3559 7500 5724 7528
rect 3559 7497 3571 7500
rect 3513 7491 3571 7497
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 5810 7488 5816 7540
rect 5868 7488 5874 7540
rect 7742 7488 7748 7540
rect 7800 7528 7806 7540
rect 7837 7531 7895 7537
rect 7837 7528 7849 7531
rect 7800 7500 7849 7528
rect 7800 7488 7806 7500
rect 7837 7497 7849 7500
rect 7883 7497 7895 7531
rect 7837 7491 7895 7497
rect 7926 7488 7932 7540
rect 7984 7528 7990 7540
rect 8113 7531 8171 7537
rect 8113 7528 8125 7531
rect 7984 7500 8125 7528
rect 7984 7488 7990 7500
rect 8113 7497 8125 7500
rect 8159 7497 8171 7531
rect 8113 7491 8171 7497
rect 4430 7460 4436 7472
rect 3068 7432 4016 7460
rect 3068 7404 3096 7432
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7392 2651 7395
rect 2869 7395 2927 7401
rect 2869 7392 2881 7395
rect 2639 7364 2881 7392
rect 2639 7361 2651 7364
rect 2593 7355 2651 7361
rect 2869 7361 2881 7364
rect 2915 7361 2927 7395
rect 2869 7355 2927 7361
rect 2961 7395 3019 7401
rect 2961 7361 2973 7395
rect 3007 7392 3019 7395
rect 3050 7392 3056 7404
rect 3007 7364 3056 7392
rect 3007 7361 3019 7364
rect 2961 7355 3019 7361
rect 3050 7352 3056 7364
rect 3108 7352 3114 7404
rect 3145 7395 3203 7401
rect 3145 7361 3157 7395
rect 3191 7392 3203 7395
rect 3234 7392 3240 7404
rect 3191 7364 3240 7392
rect 3191 7361 3203 7364
rect 3145 7355 3203 7361
rect 2317 7327 2375 7333
rect 2317 7293 2329 7327
rect 2363 7324 2375 7327
rect 3160 7324 3188 7355
rect 3234 7352 3240 7364
rect 3292 7352 3298 7404
rect 2363 7296 3188 7324
rect 2363 7293 2375 7296
rect 2317 7287 2375 7293
rect 3602 7284 3608 7336
rect 3660 7324 3666 7336
rect 3789 7327 3847 7333
rect 3789 7324 3801 7327
rect 3660 7296 3801 7324
rect 3660 7284 3666 7296
rect 3789 7293 3801 7296
rect 3835 7324 3847 7327
rect 3878 7324 3884 7336
rect 3835 7296 3884 7324
rect 3835 7293 3847 7296
rect 3789 7287 3847 7293
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 3988 7324 4016 7432
rect 4172 7432 4436 7460
rect 4065 7395 4123 7401
rect 4065 7361 4077 7395
rect 4111 7390 4123 7395
rect 4172 7390 4200 7432
rect 4430 7420 4436 7432
rect 4488 7420 4494 7472
rect 4522 7420 4528 7472
rect 4580 7420 4586 7472
rect 5828 7460 5856 7488
rect 5644 7432 5856 7460
rect 4111 7362 4200 7390
rect 4111 7361 4123 7362
rect 4065 7355 4123 7361
rect 4338 7352 4344 7404
rect 4396 7352 4402 7404
rect 4540 7333 4568 7420
rect 4617 7395 4675 7401
rect 4617 7361 4629 7395
rect 4663 7361 4675 7395
rect 4617 7355 4675 7361
rect 5445 7395 5503 7401
rect 5445 7361 5457 7395
rect 5491 7392 5503 7395
rect 5644 7392 5672 7432
rect 5491 7364 5672 7392
rect 5721 7395 5779 7401
rect 5491 7361 5503 7364
rect 5445 7355 5503 7361
rect 5721 7361 5733 7395
rect 5767 7392 5779 7395
rect 5902 7392 5908 7404
rect 5767 7364 5908 7392
rect 5767 7361 5779 7364
rect 5721 7355 5779 7361
rect 4433 7327 4491 7333
rect 3988 7296 4200 7324
rect 2501 7259 2559 7265
rect 2501 7225 2513 7259
rect 2547 7256 2559 7259
rect 3053 7259 3111 7265
rect 3053 7256 3065 7259
rect 2547 7228 3065 7256
rect 2547 7225 2559 7228
rect 2501 7219 2559 7225
rect 3053 7225 3065 7228
rect 3099 7256 3111 7259
rect 3418 7256 3424 7268
rect 3099 7228 3424 7256
rect 3099 7225 3111 7228
rect 3053 7219 3111 7225
rect 3418 7216 3424 7228
rect 3476 7216 3482 7268
rect 4062 7256 4068 7268
rect 3896 7228 4068 7256
rect 3326 7148 3332 7200
rect 3384 7188 3390 7200
rect 3896 7188 3924 7228
rect 4062 7216 4068 7228
rect 4120 7216 4126 7268
rect 4172 7256 4200 7296
rect 4433 7293 4445 7327
rect 4479 7293 4491 7327
rect 4433 7287 4491 7293
rect 4525 7327 4583 7333
rect 4525 7293 4537 7327
rect 4571 7293 4583 7327
rect 4632 7324 4660 7355
rect 5902 7352 5908 7364
rect 5960 7352 5966 7404
rect 5994 7352 6000 7404
rect 6052 7352 6058 7404
rect 6362 7352 6368 7404
rect 6420 7352 6426 7404
rect 6621 7395 6679 7401
rect 6621 7392 6633 7395
rect 6472 7364 6633 7392
rect 5626 7324 5632 7336
rect 4632 7296 5632 7324
rect 4525 7287 4583 7293
rect 4448 7256 4476 7287
rect 5626 7284 5632 7296
rect 5684 7324 5690 7336
rect 5813 7327 5871 7333
rect 5813 7324 5825 7327
rect 5684 7296 5825 7324
rect 5684 7284 5690 7296
rect 5813 7293 5825 7296
rect 5859 7293 5871 7327
rect 6472 7324 6500 7364
rect 6621 7361 6633 7364
rect 6667 7361 6679 7395
rect 6621 7355 6679 7361
rect 7374 7352 7380 7404
rect 7432 7392 7438 7404
rect 8021 7395 8079 7401
rect 8021 7392 8033 7395
rect 7432 7364 8033 7392
rect 7432 7352 7438 7364
rect 8021 7361 8033 7364
rect 8067 7361 8079 7395
rect 8021 7355 8079 7361
rect 8205 7395 8263 7401
rect 8205 7361 8217 7395
rect 8251 7361 8263 7395
rect 8205 7355 8263 7361
rect 8220 7324 8248 7355
rect 5813 7287 5871 7293
rect 6104 7296 6500 7324
rect 7760 7296 8248 7324
rect 6104 7256 6132 7296
rect 4172 7228 6132 7256
rect 3384 7160 3924 7188
rect 3973 7191 4031 7197
rect 3384 7148 3390 7160
rect 3973 7157 3985 7191
rect 4019 7188 4031 7191
rect 4157 7191 4215 7197
rect 4157 7188 4169 7191
rect 4019 7160 4169 7188
rect 4019 7157 4031 7160
rect 3973 7151 4031 7157
rect 4157 7157 4169 7160
rect 4203 7157 4215 7191
rect 4157 7151 4215 7157
rect 4338 7148 4344 7200
rect 4396 7188 4402 7200
rect 4801 7191 4859 7197
rect 4801 7188 4813 7191
rect 4396 7160 4813 7188
rect 4396 7148 4402 7160
rect 4801 7157 4813 7160
rect 4847 7157 4859 7191
rect 4801 7151 4859 7157
rect 5442 7148 5448 7200
rect 5500 7188 5506 7200
rect 5537 7191 5595 7197
rect 5537 7188 5549 7191
rect 5500 7160 5549 7188
rect 5500 7148 5506 7160
rect 5537 7157 5549 7160
rect 5583 7157 5595 7191
rect 5537 7151 5595 7157
rect 5626 7148 5632 7200
rect 5684 7188 5690 7200
rect 5736 7197 5764 7228
rect 7760 7200 7788 7296
rect 8386 7216 8392 7268
rect 8444 7216 8450 7268
rect 5721 7191 5779 7197
rect 5721 7188 5733 7191
rect 5684 7160 5733 7188
rect 5684 7148 5690 7160
rect 5721 7157 5733 7160
rect 5767 7157 5779 7191
rect 5721 7151 5779 7157
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 5994 7188 6000 7200
rect 5868 7160 6000 7188
rect 5868 7148 5874 7160
rect 5994 7148 6000 7160
rect 6052 7148 6058 7200
rect 7742 7148 7748 7200
rect 7800 7148 7806 7200
rect 1104 7098 9200 7120
rect 1104 7046 1962 7098
rect 2014 7046 2026 7098
rect 2078 7046 2090 7098
rect 2142 7046 2154 7098
rect 2206 7046 2218 7098
rect 2270 7046 3986 7098
rect 4038 7046 4050 7098
rect 4102 7046 4114 7098
rect 4166 7046 4178 7098
rect 4230 7046 4242 7098
rect 4294 7046 6010 7098
rect 6062 7046 6074 7098
rect 6126 7046 6138 7098
rect 6190 7046 6202 7098
rect 6254 7046 6266 7098
rect 6318 7046 8034 7098
rect 8086 7046 8098 7098
rect 8150 7046 8162 7098
rect 8214 7046 8226 7098
rect 8278 7046 8290 7098
rect 8342 7046 9200 7098
rect 1104 7024 9200 7046
rect 3694 6944 3700 6996
rect 3752 6984 3758 6996
rect 4065 6987 4123 6993
rect 4065 6984 4077 6987
rect 3752 6956 4077 6984
rect 3752 6944 3758 6956
rect 4065 6953 4077 6956
rect 4111 6953 4123 6987
rect 4065 6947 4123 6953
rect 5442 6944 5448 6996
rect 5500 6944 5506 6996
rect 8478 6944 8484 6996
rect 8536 6944 8542 6996
rect 5350 6916 5356 6928
rect 3528 6888 5356 6916
rect 2869 6783 2927 6789
rect 2869 6749 2881 6783
rect 2915 6780 2927 6783
rect 3326 6780 3332 6792
rect 2915 6752 3332 6780
rect 2915 6749 2927 6752
rect 2869 6743 2927 6749
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 3418 6740 3424 6792
rect 3476 6740 3482 6792
rect 3528 6780 3556 6888
rect 5350 6876 5356 6888
rect 5408 6876 5414 6928
rect 4430 6848 4436 6860
rect 4264 6820 4436 6848
rect 3602 6780 3608 6792
rect 3528 6752 3608 6780
rect 3602 6740 3608 6752
rect 3660 6740 3666 6792
rect 3694 6740 3700 6792
rect 3752 6780 3758 6792
rect 3789 6783 3847 6789
rect 3789 6780 3801 6783
rect 3752 6752 3801 6780
rect 3752 6740 3758 6752
rect 3789 6749 3801 6752
rect 3835 6780 3847 6783
rect 3878 6780 3884 6792
rect 3835 6752 3884 6780
rect 3835 6749 3847 6752
rect 3789 6743 3847 6749
rect 3878 6740 3884 6752
rect 3936 6780 3942 6792
rect 4062 6780 4068 6792
rect 3936 6752 4068 6780
rect 3936 6740 3942 6752
rect 4062 6740 4068 6752
rect 4120 6740 4126 6792
rect 4264 6789 4292 6820
rect 4430 6808 4436 6820
rect 4488 6848 4494 6860
rect 5460 6848 5488 6944
rect 7466 6876 7472 6928
rect 7524 6876 7530 6928
rect 8496 6916 8524 6944
rect 8312 6888 8524 6916
rect 4488 6820 5488 6848
rect 7837 6851 7895 6857
rect 4488 6808 4494 6820
rect 7837 6817 7849 6851
rect 7883 6848 7895 6851
rect 8113 6851 8171 6857
rect 7883 6820 8064 6848
rect 7883 6817 7895 6820
rect 7837 6811 7895 6817
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 4338 6740 4344 6792
rect 4396 6740 4402 6792
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 4617 6783 4675 6789
rect 4617 6749 4629 6783
rect 4663 6780 4675 6783
rect 5537 6783 5595 6789
rect 4663 6752 5028 6780
rect 4663 6749 4675 6752
rect 4617 6743 4675 6749
rect 2498 6672 2504 6724
rect 2556 6712 2562 6724
rect 2602 6715 2660 6721
rect 2602 6712 2614 6715
rect 2556 6684 2614 6712
rect 2556 6672 2562 6684
rect 2602 6681 2614 6684
rect 2648 6681 2660 6715
rect 2602 6675 2660 6681
rect 3513 6715 3571 6721
rect 3513 6681 3525 6715
rect 3559 6712 3571 6715
rect 4540 6712 4568 6743
rect 3559 6684 4568 6712
rect 3559 6681 3571 6684
rect 3513 6675 3571 6681
rect 5000 6656 5028 6752
rect 5537 6749 5549 6783
rect 5583 6780 5595 6783
rect 6362 6780 6368 6792
rect 5583 6752 6368 6780
rect 5583 6749 5595 6752
rect 5537 6743 5595 6749
rect 6362 6740 6368 6752
rect 6420 6740 6426 6792
rect 7193 6783 7251 6789
rect 7193 6749 7205 6783
rect 7239 6780 7251 6783
rect 7745 6783 7803 6789
rect 7239 6752 7420 6780
rect 7239 6749 7251 6752
rect 7193 6743 7251 6749
rect 7392 6724 7420 6752
rect 7745 6749 7757 6783
rect 7791 6780 7803 6783
rect 7926 6780 7932 6792
rect 7791 6752 7932 6780
rect 7791 6749 7803 6752
rect 7745 6743 7803 6749
rect 7926 6740 7932 6752
rect 7984 6740 7990 6792
rect 8036 6780 8064 6820
rect 8113 6817 8125 6851
rect 8159 6848 8171 6851
rect 8312 6848 8340 6888
rect 8159 6820 8340 6848
rect 8389 6851 8447 6857
rect 8159 6817 8171 6820
rect 8113 6811 8171 6817
rect 8389 6817 8401 6851
rect 8435 6848 8447 6851
rect 8570 6848 8576 6860
rect 8435 6820 8576 6848
rect 8435 6817 8447 6820
rect 8389 6811 8447 6817
rect 8570 6808 8576 6820
rect 8628 6808 8634 6860
rect 8478 6780 8484 6792
rect 8036 6752 8484 6780
rect 8478 6740 8484 6752
rect 8536 6740 8542 6792
rect 5804 6715 5862 6721
rect 5804 6681 5816 6715
rect 5850 6712 5862 6715
rect 5902 6712 5908 6724
rect 5850 6684 5908 6712
rect 5850 6681 5862 6684
rect 5804 6675 5862 6681
rect 5902 6672 5908 6684
rect 5960 6672 5966 6724
rect 7374 6672 7380 6724
rect 7432 6672 7438 6724
rect 7469 6715 7527 6721
rect 7469 6681 7481 6715
rect 7515 6712 7527 6715
rect 7650 6712 7656 6724
rect 7515 6684 7656 6712
rect 7515 6681 7527 6684
rect 7469 6675 7527 6681
rect 7650 6672 7656 6684
rect 7708 6672 7714 6724
rect 8665 6715 8723 6721
rect 8665 6681 8677 6715
rect 8711 6712 8723 6715
rect 8711 6684 9260 6712
rect 8711 6681 8723 6684
rect 8665 6675 8723 6681
rect 1486 6604 1492 6656
rect 1544 6604 1550 6656
rect 3050 6604 3056 6656
rect 3108 6644 3114 6656
rect 3694 6644 3700 6656
rect 3108 6616 3700 6644
rect 3108 6604 3114 6616
rect 3694 6604 3700 6616
rect 3752 6604 3758 6656
rect 3878 6604 3884 6656
rect 3936 6604 3942 6656
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 4982 6644 4988 6656
rect 4120 6616 4988 6644
rect 4120 6604 4126 6616
rect 4982 6604 4988 6616
rect 5040 6604 5046 6656
rect 6917 6647 6975 6653
rect 6917 6613 6929 6647
rect 6963 6644 6975 6647
rect 7285 6647 7343 6653
rect 7285 6644 7297 6647
rect 6963 6616 7297 6644
rect 6963 6613 6975 6616
rect 6917 6607 6975 6613
rect 7285 6613 7297 6616
rect 7331 6644 7343 6647
rect 8386 6644 8392 6656
rect 7331 6616 8392 6644
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 1104 6554 9200 6576
rect 1104 6502 2622 6554
rect 2674 6502 2686 6554
rect 2738 6502 2750 6554
rect 2802 6502 2814 6554
rect 2866 6502 2878 6554
rect 2930 6502 4646 6554
rect 4698 6502 4710 6554
rect 4762 6502 4774 6554
rect 4826 6502 4838 6554
rect 4890 6502 4902 6554
rect 4954 6502 6670 6554
rect 6722 6502 6734 6554
rect 6786 6502 6798 6554
rect 6850 6502 6862 6554
rect 6914 6502 6926 6554
rect 6978 6502 8694 6554
rect 8746 6502 8758 6554
rect 8810 6502 8822 6554
rect 8874 6502 8886 6554
rect 8938 6502 8950 6554
rect 9002 6502 9200 6554
rect 1104 6480 9200 6502
rect 1486 6400 1492 6452
rect 1544 6400 1550 6452
rect 3326 6400 3332 6452
rect 3384 6440 3390 6452
rect 3384 6412 3832 6440
rect 3384 6400 3390 6412
rect 1504 6304 1532 6400
rect 1765 6307 1823 6313
rect 1765 6304 1777 6307
rect 1504 6276 1777 6304
rect 1765 6273 1777 6276
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 2961 6307 3019 6313
rect 2961 6273 2973 6307
rect 3007 6304 3019 6307
rect 3234 6304 3240 6316
rect 3007 6276 3240 6304
rect 3007 6273 3019 6276
rect 2961 6267 3019 6273
rect 3234 6264 3240 6276
rect 3292 6264 3298 6316
rect 3421 6307 3479 6313
rect 3421 6273 3433 6307
rect 3467 6273 3479 6307
rect 3421 6267 3479 6273
rect 3436 6236 3464 6267
rect 3602 6264 3608 6316
rect 3660 6264 3666 6316
rect 3620 6236 3648 6264
rect 2424 6208 3464 6236
rect 3528 6208 3648 6236
rect 3804 6236 3832 6412
rect 5166 6400 5172 6452
rect 5224 6440 5230 6452
rect 5997 6443 6055 6449
rect 5997 6440 6009 6443
rect 5224 6412 6009 6440
rect 5224 6400 5230 6412
rect 5997 6409 6009 6412
rect 6043 6409 6055 6443
rect 5997 6403 6055 6409
rect 7466 6400 7472 6452
rect 7524 6440 7530 6452
rect 8757 6443 8815 6449
rect 7524 6412 8708 6440
rect 7524 6400 7530 6412
rect 4062 6332 4068 6384
rect 4120 6372 4126 6384
rect 8205 6375 8263 6381
rect 8205 6372 8217 6375
rect 4120 6344 5856 6372
rect 4120 6332 4126 6344
rect 3973 6307 4031 6313
rect 3973 6273 3985 6307
rect 4019 6304 4031 6307
rect 4080 6304 4108 6332
rect 5828 6316 5856 6344
rect 7944 6344 8217 6372
rect 4338 6313 4344 6316
rect 4019 6276 4108 6304
rect 4019 6273 4031 6276
rect 3973 6267 4031 6273
rect 4332 6267 4344 6313
rect 4338 6264 4344 6267
rect 4396 6264 4402 6316
rect 5810 6264 5816 6316
rect 5868 6264 5874 6316
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6273 6239 6307
rect 6181 6267 6239 6273
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6304 7619 6307
rect 7944 6304 7972 6344
rect 8205 6341 8217 6344
rect 8251 6372 8263 6375
rect 8294 6372 8300 6384
rect 8251 6344 8300 6372
rect 8251 6341 8263 6344
rect 8205 6335 8263 6341
rect 8294 6332 8300 6344
rect 8352 6332 8358 6384
rect 8405 6375 8463 6381
rect 8405 6372 8417 6375
rect 8404 6341 8417 6372
rect 8451 6341 8463 6375
rect 8404 6335 8463 6341
rect 7607 6276 7972 6304
rect 7607 6273 7619 6276
rect 7561 6267 7619 6273
rect 4065 6239 4123 6245
rect 4065 6236 4077 6239
rect 3804 6208 4077 6236
rect 2424 6112 2452 6208
rect 3142 6128 3148 6180
rect 3200 6168 3206 6180
rect 3528 6168 3556 6208
rect 4065 6205 4077 6208
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 3200 6140 3556 6168
rect 3200 6128 3206 6140
rect 3602 6128 3608 6180
rect 3660 6168 3666 6180
rect 5445 6171 5503 6177
rect 3660 6140 3924 6168
rect 3660 6128 3666 6140
rect 2406 6060 2412 6112
rect 2464 6060 2470 6112
rect 2682 6060 2688 6112
rect 2740 6060 2746 6112
rect 3050 6060 3056 6112
rect 3108 6060 3114 6112
rect 3237 6103 3295 6109
rect 3237 6069 3249 6103
rect 3283 6100 3295 6103
rect 3418 6100 3424 6112
rect 3283 6072 3424 6100
rect 3283 6069 3295 6072
rect 3237 6063 3295 6069
rect 3418 6060 3424 6072
rect 3476 6100 3482 6112
rect 3789 6103 3847 6109
rect 3789 6100 3801 6103
rect 3476 6072 3801 6100
rect 3476 6060 3482 6072
rect 3789 6069 3801 6072
rect 3835 6069 3847 6103
rect 3896 6100 3924 6140
rect 5445 6137 5457 6171
rect 5491 6168 5503 6171
rect 6196 6168 6224 6267
rect 7374 6196 7380 6248
rect 7432 6236 7438 6248
rect 7653 6239 7711 6245
rect 7653 6236 7665 6239
rect 7432 6208 7665 6236
rect 7432 6196 7438 6208
rect 7653 6205 7665 6208
rect 7699 6236 7711 6239
rect 8404 6236 8432 6335
rect 8680 6313 8708 6412
rect 8757 6409 8769 6443
rect 8803 6440 8815 6443
rect 9232 6440 9260 6684
rect 8803 6412 9260 6440
rect 8803 6409 8815 6412
rect 8757 6403 8815 6409
rect 8665 6307 8723 6313
rect 8665 6273 8677 6307
rect 8711 6273 8723 6307
rect 8665 6267 8723 6273
rect 8849 6307 8907 6313
rect 8849 6273 8861 6307
rect 8895 6273 8907 6307
rect 8849 6267 8907 6273
rect 7699 6208 8432 6236
rect 7699 6205 7711 6208
rect 7653 6199 7711 6205
rect 5491 6140 6224 6168
rect 5491 6137 5503 6140
rect 5445 6131 5503 6137
rect 4062 6100 4068 6112
rect 3896 6072 4068 6100
rect 3789 6063 3847 6069
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 4430 6060 4436 6112
rect 4488 6100 4494 6112
rect 5460 6100 5488 6131
rect 4488 6072 5488 6100
rect 7668 6100 7696 6199
rect 8478 6196 8484 6248
rect 8536 6236 8542 6248
rect 8864 6236 8892 6267
rect 8536 6208 8892 6236
rect 8536 6196 8542 6208
rect 8496 6168 8524 6196
rect 8573 6171 8631 6177
rect 8573 6168 8585 6171
rect 8496 6140 8585 6168
rect 8573 6137 8585 6140
rect 8619 6137 8631 6171
rect 8573 6131 8631 6137
rect 7834 6100 7840 6112
rect 7668 6072 7840 6100
rect 4488 6060 4494 6072
rect 7834 6060 7840 6072
rect 7892 6060 7898 6112
rect 7926 6060 7932 6112
rect 7984 6060 7990 6112
rect 8018 6060 8024 6112
rect 8076 6100 8082 6112
rect 8389 6103 8447 6109
rect 8389 6100 8401 6103
rect 8076 6072 8401 6100
rect 8076 6060 8082 6072
rect 8389 6069 8401 6072
rect 8435 6069 8447 6103
rect 8389 6063 8447 6069
rect 1104 6010 9200 6032
rect 1104 5958 1962 6010
rect 2014 5958 2026 6010
rect 2078 5958 2090 6010
rect 2142 5958 2154 6010
rect 2206 5958 2218 6010
rect 2270 5958 3986 6010
rect 4038 5958 4050 6010
rect 4102 5958 4114 6010
rect 4166 5958 4178 6010
rect 4230 5958 4242 6010
rect 4294 5958 6010 6010
rect 6062 5958 6074 6010
rect 6126 5958 6138 6010
rect 6190 5958 6202 6010
rect 6254 5958 6266 6010
rect 6318 5958 8034 6010
rect 8086 5958 8098 6010
rect 8150 5958 8162 6010
rect 8214 5958 8226 6010
rect 8278 5958 8290 6010
rect 8342 5958 9200 6010
rect 1104 5936 9200 5958
rect 750 5856 756 5908
rect 808 5896 814 5908
rect 1489 5899 1547 5905
rect 1489 5896 1501 5899
rect 808 5868 1501 5896
rect 808 5856 814 5868
rect 1489 5865 1501 5868
rect 1535 5865 1547 5899
rect 1489 5859 1547 5865
rect 2409 5899 2467 5905
rect 2409 5865 2421 5899
rect 2455 5896 2467 5899
rect 2498 5896 2504 5908
rect 2455 5868 2504 5896
rect 2455 5865 2467 5868
rect 2409 5859 2467 5865
rect 2498 5856 2504 5868
rect 2556 5856 2562 5908
rect 2682 5856 2688 5908
rect 2740 5856 2746 5908
rect 3142 5896 3148 5908
rect 2792 5868 3148 5896
rect 1486 5720 1492 5772
rect 1544 5720 1550 5772
rect 2406 5760 2412 5772
rect 2148 5732 2412 5760
rect 1504 5692 1532 5720
rect 2148 5701 2176 5732
rect 2406 5720 2412 5732
rect 2464 5720 2470 5772
rect 2501 5763 2559 5769
rect 2501 5729 2513 5763
rect 2547 5760 2559 5763
rect 2700 5760 2728 5856
rect 2792 5837 2820 5868
rect 3142 5856 3148 5868
rect 3200 5856 3206 5908
rect 3234 5856 3240 5908
rect 3292 5896 3298 5908
rect 3878 5896 3884 5908
rect 3292 5868 3884 5896
rect 3292 5856 3298 5868
rect 3878 5856 3884 5868
rect 3936 5856 3942 5908
rect 5074 5856 5080 5908
rect 5132 5856 5138 5908
rect 7926 5856 7932 5908
rect 7984 5856 7990 5908
rect 8662 5856 8668 5908
rect 8720 5856 8726 5908
rect 2777 5831 2835 5837
rect 2777 5797 2789 5831
rect 2823 5797 2835 5831
rect 2777 5791 2835 5797
rect 3418 5760 3424 5772
rect 2547 5732 2728 5760
rect 2792 5732 3424 5760
rect 2547 5729 2559 5732
rect 2501 5723 2559 5729
rect 1765 5695 1823 5701
rect 1765 5692 1777 5695
rect 1504 5664 1777 5692
rect 1765 5661 1777 5664
rect 1811 5661 1823 5695
rect 1765 5655 1823 5661
rect 2133 5695 2191 5701
rect 2133 5661 2145 5695
rect 2179 5661 2191 5695
rect 2133 5655 2191 5661
rect 2225 5695 2283 5701
rect 2225 5661 2237 5695
rect 2271 5661 2283 5695
rect 2225 5655 2283 5661
rect 2317 5695 2375 5701
rect 2317 5661 2329 5695
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 2593 5695 2651 5701
rect 2593 5661 2605 5695
rect 2639 5692 2651 5695
rect 2792 5692 2820 5732
rect 3418 5720 3424 5732
rect 3476 5720 3482 5772
rect 2639 5664 2820 5692
rect 2869 5695 2927 5701
rect 2639 5661 2651 5664
rect 2593 5655 2651 5661
rect 2869 5661 2881 5695
rect 2915 5692 2927 5695
rect 3050 5692 3056 5704
rect 2915 5664 3056 5692
rect 2915 5661 2927 5664
rect 2869 5655 2927 5661
rect 2041 5627 2099 5633
rect 2041 5593 2053 5627
rect 2087 5624 2099 5627
rect 2240 5624 2268 5655
rect 2087 5596 2268 5624
rect 2087 5593 2099 5596
rect 2041 5587 2099 5593
rect 2332 5556 2360 5655
rect 3050 5652 3056 5664
rect 3108 5692 3114 5704
rect 3108 5664 3740 5692
rect 3108 5652 3114 5664
rect 3712 5636 3740 5664
rect 3786 5652 3792 5704
rect 3844 5652 3850 5704
rect 6178 5652 6184 5704
rect 6236 5652 6242 5704
rect 7650 5652 7656 5704
rect 7708 5652 7714 5704
rect 7837 5695 7895 5701
rect 7837 5661 7849 5695
rect 7883 5661 7895 5695
rect 7944 5692 7972 5856
rect 8481 5695 8539 5701
rect 8481 5692 8493 5695
rect 7944 5664 8493 5692
rect 7837 5655 7895 5661
rect 8481 5661 8493 5664
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 3694 5584 3700 5636
rect 3752 5584 3758 5636
rect 7852 5624 7880 5655
rect 7926 5624 7932 5636
rect 7852 5596 7932 5624
rect 7926 5584 7932 5596
rect 7984 5584 7990 5636
rect 2406 5556 2412 5568
rect 2332 5528 2412 5556
rect 2406 5516 2412 5528
rect 2464 5556 2470 5568
rect 2869 5559 2927 5565
rect 2869 5556 2881 5559
rect 2464 5528 2881 5556
rect 2464 5516 2470 5528
rect 2869 5525 2881 5528
rect 2915 5525 2927 5559
rect 2869 5519 2927 5525
rect 5626 5516 5632 5568
rect 5684 5516 5690 5568
rect 7745 5559 7803 5565
rect 7745 5525 7757 5559
rect 7791 5556 7803 5559
rect 8294 5556 8300 5568
rect 7791 5528 8300 5556
rect 7791 5525 7803 5528
rect 7745 5519 7803 5525
rect 8294 5516 8300 5528
rect 8352 5516 8358 5568
rect 1104 5466 9200 5488
rect 1104 5414 2622 5466
rect 2674 5414 2686 5466
rect 2738 5414 2750 5466
rect 2802 5414 2814 5466
rect 2866 5414 2878 5466
rect 2930 5414 4646 5466
rect 4698 5414 4710 5466
rect 4762 5414 4774 5466
rect 4826 5414 4838 5466
rect 4890 5414 4902 5466
rect 4954 5414 6670 5466
rect 6722 5414 6734 5466
rect 6786 5414 6798 5466
rect 6850 5414 6862 5466
rect 6914 5414 6926 5466
rect 6978 5414 8694 5466
rect 8746 5414 8758 5466
rect 8810 5414 8822 5466
rect 8874 5414 8886 5466
rect 8938 5414 8950 5466
rect 9002 5414 9200 5466
rect 1104 5392 9200 5414
rect 3694 5312 3700 5364
rect 3752 5312 3758 5364
rect 4065 5355 4123 5361
rect 4065 5321 4077 5355
rect 4111 5352 4123 5355
rect 4338 5352 4344 5364
rect 4111 5324 4344 5352
rect 4111 5321 4123 5324
rect 4065 5315 4123 5321
rect 4338 5312 4344 5324
rect 4396 5312 4402 5364
rect 5166 5312 5172 5364
rect 5224 5312 5230 5364
rect 3050 5284 3056 5296
rect 2148 5256 3056 5284
rect 2148 5225 2176 5256
rect 3050 5244 3056 5256
rect 3108 5244 3114 5296
rect 5184 5284 5212 5312
rect 4172 5256 5212 5284
rect 2133 5219 2191 5225
rect 2133 5185 2145 5219
rect 2179 5185 2191 5219
rect 2133 5179 2191 5185
rect 2225 5219 2283 5225
rect 2225 5185 2237 5219
rect 2271 5185 2283 5219
rect 2225 5179 2283 5185
rect 2240 5148 2268 5179
rect 2406 5176 2412 5228
rect 2464 5176 2470 5228
rect 2498 5176 2504 5228
rect 2556 5176 2562 5228
rect 3329 5219 3387 5225
rect 3329 5216 3341 5219
rect 3160 5188 3341 5216
rect 3160 5157 3188 5188
rect 3329 5185 3341 5188
rect 3375 5185 3387 5219
rect 3329 5179 3387 5185
rect 3510 5176 3516 5228
rect 3568 5176 3574 5228
rect 3878 5176 3884 5228
rect 3936 5216 3942 5228
rect 4172 5225 4200 5256
rect 3973 5219 4031 5225
rect 3973 5216 3985 5219
rect 3936 5188 3985 5216
rect 3936 5176 3942 5188
rect 3973 5185 3985 5188
rect 4019 5185 4031 5219
rect 3973 5179 4031 5185
rect 4157 5219 4215 5225
rect 4157 5185 4169 5219
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 4700 5219 4758 5225
rect 4700 5185 4712 5219
rect 4746 5216 4758 5219
rect 5166 5216 5172 5228
rect 4746 5188 5172 5216
rect 4746 5185 4758 5188
rect 4700 5179 4758 5185
rect 5166 5176 5172 5188
rect 5224 5176 5230 5228
rect 6178 5216 6184 5228
rect 5828 5188 6184 5216
rect 2593 5151 2651 5157
rect 2593 5148 2605 5151
rect 2240 5120 2605 5148
rect 2593 5117 2605 5120
rect 2639 5117 2651 5151
rect 3145 5151 3203 5157
rect 3145 5148 3157 5151
rect 2593 5111 2651 5117
rect 2792 5120 3157 5148
rect 2792 5024 2820 5120
rect 3145 5117 3157 5120
rect 3191 5117 3203 5151
rect 3145 5111 3203 5117
rect 4430 5108 4436 5160
rect 4488 5108 4494 5160
rect 1670 4972 1676 5024
rect 1728 5012 1734 5024
rect 1949 5015 2007 5021
rect 1949 5012 1961 5015
rect 1728 4984 1961 5012
rect 1728 4972 1734 4984
rect 1949 4981 1961 4984
rect 1995 4981 2007 5015
rect 1949 4975 2007 4981
rect 2774 4972 2780 5024
rect 2832 4972 2838 5024
rect 4706 4972 4712 5024
rect 4764 5012 4770 5024
rect 5828 5021 5856 5188
rect 6178 5176 6184 5188
rect 6236 5216 6242 5228
rect 6621 5219 6679 5225
rect 6621 5216 6633 5219
rect 6236 5188 6633 5216
rect 6236 5176 6242 5188
rect 6621 5185 6633 5188
rect 6667 5185 6679 5219
rect 6621 5179 6679 5185
rect 7466 5176 7472 5228
rect 7524 5216 7530 5228
rect 8021 5219 8079 5225
rect 8021 5216 8033 5219
rect 7524 5188 8033 5216
rect 7524 5176 7530 5188
rect 8021 5185 8033 5188
rect 8067 5185 8079 5219
rect 8021 5179 8079 5185
rect 8294 5176 8300 5228
rect 8352 5216 8358 5228
rect 8573 5219 8631 5225
rect 8573 5216 8585 5219
rect 8352 5188 8585 5216
rect 8352 5176 8358 5188
rect 8573 5185 8585 5188
rect 8619 5185 8631 5219
rect 8573 5179 8631 5185
rect 6362 5108 6368 5160
rect 6420 5108 6426 5160
rect 7834 5108 7840 5160
rect 7892 5148 7898 5160
rect 7929 5151 7987 5157
rect 7929 5148 7941 5151
rect 7892 5120 7941 5148
rect 7892 5108 7898 5120
rect 7929 5117 7941 5120
rect 7975 5117 7987 5151
rect 7929 5111 7987 5117
rect 5813 5015 5871 5021
rect 5813 5012 5825 5015
rect 4764 4984 5825 5012
rect 4764 4972 4770 4984
rect 5813 4981 5825 4984
rect 5859 4981 5871 5015
rect 5813 4975 5871 4981
rect 7742 4972 7748 5024
rect 7800 4972 7806 5024
rect 8297 5015 8355 5021
rect 8297 4981 8309 5015
rect 8343 5012 8355 5015
rect 8386 5012 8392 5024
rect 8343 4984 8392 5012
rect 8343 4981 8355 4984
rect 8297 4975 8355 4981
rect 8386 4972 8392 4984
rect 8444 4972 8450 5024
rect 8754 4972 8760 5024
rect 8812 4972 8818 5024
rect 1104 4922 9200 4944
rect 1104 4870 1962 4922
rect 2014 4870 2026 4922
rect 2078 4870 2090 4922
rect 2142 4870 2154 4922
rect 2206 4870 2218 4922
rect 2270 4870 3986 4922
rect 4038 4870 4050 4922
rect 4102 4870 4114 4922
rect 4166 4870 4178 4922
rect 4230 4870 4242 4922
rect 4294 4870 6010 4922
rect 6062 4870 6074 4922
rect 6126 4870 6138 4922
rect 6190 4870 6202 4922
rect 6254 4870 6266 4922
rect 6318 4870 8034 4922
rect 8086 4870 8098 4922
rect 8150 4870 8162 4922
rect 8214 4870 8226 4922
rect 8278 4870 8290 4922
rect 8342 4870 9200 4922
rect 1104 4848 9200 4870
rect 2774 4768 2780 4820
rect 2832 4768 2838 4820
rect 3142 4808 3148 4820
rect 2976 4780 3148 4808
rect 1394 4564 1400 4616
rect 1452 4564 1458 4616
rect 1670 4613 1676 4616
rect 1664 4604 1676 4613
rect 1631 4576 1676 4604
rect 1664 4567 1676 4576
rect 1670 4564 1676 4567
rect 1728 4564 1734 4616
rect 2976 4536 3004 4780
rect 3142 4768 3148 4780
rect 3200 4808 3206 4820
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 3200 4780 3249 4808
rect 3200 4768 3206 4780
rect 3237 4777 3249 4780
rect 3283 4777 3295 4811
rect 3237 4771 3295 4777
rect 3602 4768 3608 4820
rect 3660 4808 3666 4820
rect 3973 4811 4031 4817
rect 3973 4808 3985 4811
rect 3660 4780 3985 4808
rect 3660 4768 3666 4780
rect 3973 4777 3985 4780
rect 4019 4808 4031 4811
rect 4249 4811 4307 4817
rect 4249 4808 4261 4811
rect 4019 4780 4261 4808
rect 4019 4777 4031 4780
rect 3973 4771 4031 4777
rect 4249 4777 4261 4780
rect 4295 4777 4307 4811
rect 4249 4771 4307 4777
rect 4522 4768 4528 4820
rect 4580 4768 4586 4820
rect 5166 4768 5172 4820
rect 5224 4808 5230 4820
rect 5261 4811 5319 4817
rect 5261 4808 5273 4811
rect 5224 4780 5273 4808
rect 5224 4768 5230 4780
rect 5261 4777 5273 4780
rect 5307 4777 5319 4811
rect 5261 4771 5319 4777
rect 7561 4811 7619 4817
rect 7561 4777 7573 4811
rect 7607 4808 7619 4811
rect 7650 4808 7656 4820
rect 7607 4780 7656 4808
rect 7607 4777 7619 4780
rect 7561 4771 7619 4777
rect 7650 4768 7656 4780
rect 7708 4768 7714 4820
rect 8386 4768 8392 4820
rect 8444 4768 8450 4820
rect 3050 4700 3056 4752
rect 3108 4740 3114 4752
rect 3789 4743 3847 4749
rect 3789 4740 3801 4743
rect 3108 4712 3801 4740
rect 3108 4700 3114 4712
rect 3789 4709 3801 4712
rect 3835 4709 3847 4743
rect 5077 4743 5135 4749
rect 3789 4703 3847 4709
rect 3896 4712 5028 4740
rect 3053 4607 3111 4613
rect 3053 4573 3065 4607
rect 3099 4604 3111 4607
rect 3142 4604 3148 4616
rect 3099 4576 3148 4604
rect 3099 4573 3111 4576
rect 3053 4567 3111 4573
rect 3142 4564 3148 4576
rect 3200 4564 3206 4616
rect 3329 4607 3387 4613
rect 3329 4573 3341 4607
rect 3375 4604 3387 4607
rect 3418 4604 3424 4616
rect 3375 4576 3424 4604
rect 3375 4573 3387 4576
rect 3329 4567 3387 4573
rect 3418 4564 3424 4576
rect 3476 4604 3482 4616
rect 3896 4604 3924 4712
rect 5000 4672 5028 4712
rect 5077 4709 5089 4743
rect 5123 4740 5135 4743
rect 7009 4743 7067 4749
rect 5123 4712 5304 4740
rect 5123 4709 5135 4712
rect 5077 4703 5135 4709
rect 4264 4644 4844 4672
rect 5000 4644 5212 4672
rect 3476 4576 3924 4604
rect 3476 4564 3482 4576
rect 3970 4564 3976 4616
rect 4028 4564 4034 4616
rect 4157 4607 4215 4613
rect 4157 4573 4169 4607
rect 4203 4573 4215 4607
rect 4157 4567 4215 4573
rect 4172 4536 4200 4567
rect 2976 4508 4200 4536
rect 4264 4536 4292 4644
rect 4338 4564 4344 4616
rect 4396 4604 4402 4616
rect 4433 4607 4491 4613
rect 4433 4604 4445 4607
rect 4396 4576 4445 4604
rect 4396 4564 4402 4576
rect 4433 4573 4445 4576
rect 4479 4573 4491 4607
rect 4433 4567 4491 4573
rect 4525 4607 4583 4613
rect 4525 4573 4537 4607
rect 4571 4573 4583 4607
rect 4525 4567 4583 4573
rect 4540 4536 4568 4567
rect 4706 4564 4712 4616
rect 4764 4564 4770 4616
rect 4816 4613 4844 4644
rect 4801 4607 4859 4613
rect 4801 4573 4813 4607
rect 4847 4573 4859 4607
rect 4801 4567 4859 4573
rect 4890 4564 4896 4616
rect 4948 4604 4954 4616
rect 5184 4613 5212 4644
rect 5077 4607 5135 4613
rect 5077 4604 5089 4607
rect 4948 4576 5089 4604
rect 4948 4564 4954 4576
rect 5077 4573 5089 4576
rect 5123 4573 5135 4607
rect 5077 4567 5135 4573
rect 5169 4607 5227 4613
rect 5169 4573 5181 4607
rect 5215 4573 5227 4607
rect 5276 4604 5304 4712
rect 7009 4709 7021 4743
rect 7055 4740 7067 4743
rect 7466 4740 7472 4752
rect 7055 4712 7472 4740
rect 7055 4709 7067 4712
rect 7009 4703 7067 4709
rect 5353 4607 5411 4613
rect 5353 4604 5365 4607
rect 5276 4576 5365 4604
rect 5169 4567 5227 4573
rect 5353 4573 5365 4576
rect 5399 4573 5411 4607
rect 5353 4567 5411 4573
rect 5629 4607 5687 4613
rect 5629 4573 5641 4607
rect 5675 4604 5687 4607
rect 6362 4604 6368 4616
rect 5675 4576 6368 4604
rect 5675 4573 5687 4576
rect 5629 4567 5687 4573
rect 6362 4564 6368 4576
rect 6420 4564 6426 4616
rect 7300 4613 7328 4712
rect 7466 4700 7472 4712
rect 7524 4700 7530 4752
rect 7377 4675 7435 4681
rect 7377 4641 7389 4675
rect 7423 4672 7435 4675
rect 7423 4644 8248 4672
rect 7423 4641 7435 4644
rect 7377 4635 7435 4641
rect 7285 4607 7343 4613
rect 7285 4573 7297 4607
rect 7331 4573 7343 4607
rect 7285 4567 7343 4573
rect 7742 4564 7748 4616
rect 7800 4564 7806 4616
rect 7834 4564 7840 4616
rect 7892 4604 7898 4616
rect 8220 4613 8248 4644
rect 8021 4607 8079 4613
rect 8021 4604 8033 4607
rect 7892 4576 8033 4604
rect 7892 4564 7898 4576
rect 8021 4573 8033 4576
rect 8067 4573 8079 4607
rect 8021 4567 8079 4573
rect 8205 4607 8263 4613
rect 8205 4573 8217 4607
rect 8251 4573 8263 4607
rect 8404 4604 8432 4768
rect 8481 4607 8539 4613
rect 8481 4604 8493 4607
rect 8404 4576 8493 4604
rect 8205 4567 8263 4573
rect 8481 4573 8493 4576
rect 8527 4573 8539 4607
rect 8481 4567 8539 4573
rect 4982 4536 4988 4548
rect 4264 4508 4384 4536
rect 4540 4508 4988 4536
rect 4356 4480 4384 4508
rect 4982 4496 4988 4508
rect 5040 4536 5046 4548
rect 5874 4539 5932 4545
rect 5874 4536 5886 4539
rect 5040 4508 5886 4536
rect 5040 4496 5046 4508
rect 5874 4505 5886 4508
rect 5920 4505 5932 4539
rect 5874 4499 5932 4505
rect 2869 4471 2927 4477
rect 2869 4437 2881 4471
rect 2915 4468 2927 4471
rect 2958 4468 2964 4480
rect 2915 4440 2964 4468
rect 2915 4437 2927 4440
rect 2869 4431 2927 4437
rect 2958 4428 2964 4440
rect 3016 4428 3022 4480
rect 3142 4428 3148 4480
rect 3200 4468 3206 4480
rect 3510 4468 3516 4480
rect 3200 4440 3516 4468
rect 3200 4428 3206 4440
rect 3510 4428 3516 4440
rect 3568 4468 3574 4480
rect 3970 4468 3976 4480
rect 3568 4440 3976 4468
rect 3568 4428 3574 4440
rect 3970 4428 3976 4440
rect 4028 4428 4034 4480
rect 4338 4428 4344 4480
rect 4396 4428 4402 4480
rect 4893 4471 4951 4477
rect 4893 4437 4905 4471
rect 4939 4468 4951 4471
rect 5626 4468 5632 4480
rect 4939 4440 5632 4468
rect 4939 4437 4951 4440
rect 4893 4431 4951 4437
rect 5626 4428 5632 4440
rect 5684 4428 5690 4480
rect 8665 4471 8723 4477
rect 8665 4437 8677 4471
rect 8711 4468 8723 4471
rect 9122 4468 9128 4480
rect 8711 4440 9128 4468
rect 8711 4437 8723 4440
rect 8665 4431 8723 4437
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 1104 4378 9200 4400
rect 1104 4326 2622 4378
rect 2674 4326 2686 4378
rect 2738 4326 2750 4378
rect 2802 4326 2814 4378
rect 2866 4326 2878 4378
rect 2930 4326 4646 4378
rect 4698 4326 4710 4378
rect 4762 4326 4774 4378
rect 4826 4326 4838 4378
rect 4890 4326 4902 4378
rect 4954 4326 6670 4378
rect 6722 4326 6734 4378
rect 6786 4326 6798 4378
rect 6850 4326 6862 4378
rect 6914 4326 6926 4378
rect 6978 4326 8694 4378
rect 8746 4326 8758 4378
rect 8810 4326 8822 4378
rect 8874 4326 8886 4378
rect 8938 4326 8950 4378
rect 9002 4326 9200 4378
rect 1104 4304 9200 4326
rect 3050 4224 3056 4276
rect 3108 4224 3114 4276
rect 4246 4224 4252 4276
rect 4304 4264 4310 4276
rect 4706 4264 4712 4276
rect 4304 4236 4712 4264
rect 4304 4224 4310 4236
rect 4706 4224 4712 4236
rect 4764 4224 4770 4276
rect 5166 4224 5172 4276
rect 5224 4224 5230 4276
rect 7742 4224 7748 4276
rect 7800 4224 7806 4276
rect 2777 4131 2835 4137
rect 2777 4097 2789 4131
rect 2823 4128 2835 4131
rect 3068 4128 3096 4224
rect 5184 4137 5212 4224
rect 7760 4196 7788 4224
rect 7484 4168 7788 4196
rect 7484 4137 7512 4168
rect 2823 4100 3096 4128
rect 5169 4131 5227 4137
rect 2823 4097 2835 4100
rect 2777 4091 2835 4097
rect 5169 4097 5181 4131
rect 5215 4097 5227 4131
rect 5169 4091 5227 4097
rect 7469 4131 7527 4137
rect 7469 4097 7481 4131
rect 7515 4097 7527 4131
rect 7469 4091 7527 4097
rect 7558 4088 7564 4140
rect 7616 4128 7622 4140
rect 7653 4131 7711 4137
rect 7653 4128 7665 4131
rect 7616 4100 7665 4128
rect 7616 4088 7622 4100
rect 7653 4097 7665 4100
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 7742 4088 7748 4140
rect 7800 4088 7806 4140
rect 7837 4131 7895 4137
rect 7837 4097 7849 4131
rect 7883 4097 7895 4131
rect 7837 4091 7895 4097
rect 2498 4020 2504 4072
rect 2556 4020 2562 4072
rect 4522 4020 4528 4072
rect 4580 4060 4586 4072
rect 4893 4063 4951 4069
rect 4893 4060 4905 4063
rect 4580 4032 4905 4060
rect 4580 4020 4586 4032
rect 4893 4029 4905 4032
rect 4939 4029 4951 4063
rect 7852 4060 7880 4091
rect 4893 4023 4951 4029
rect 7668 4032 7880 4060
rect 7668 3936 7696 4032
rect 7926 4020 7932 4072
rect 7984 4060 7990 4072
rect 8113 4063 8171 4069
rect 8113 4060 8125 4063
rect 7984 4032 8125 4060
rect 7984 4020 7990 4032
rect 8113 4029 8125 4032
rect 8159 4029 8171 4063
rect 8113 4023 8171 4029
rect 2225 3927 2283 3933
rect 2225 3893 2237 3927
rect 2271 3924 2283 3927
rect 2314 3924 2320 3936
rect 2271 3896 2320 3924
rect 2271 3893 2283 3896
rect 2225 3887 2283 3893
rect 2314 3884 2320 3896
rect 2372 3884 2378 3936
rect 2685 3927 2743 3933
rect 2685 3893 2697 3927
rect 2731 3924 2743 3927
rect 2958 3924 2964 3936
rect 2731 3896 2964 3924
rect 2731 3893 2743 3896
rect 2685 3887 2743 3893
rect 2958 3884 2964 3896
rect 3016 3884 3022 3936
rect 4982 3884 4988 3936
rect 5040 3884 5046 3936
rect 5077 3927 5135 3933
rect 5077 3893 5089 3927
rect 5123 3924 5135 3927
rect 5166 3924 5172 3936
rect 5123 3896 5172 3924
rect 5123 3893 5135 3896
rect 5077 3887 5135 3893
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 7650 3884 7656 3936
rect 7708 3884 7714 3936
rect 1104 3834 9200 3856
rect 1104 3782 1962 3834
rect 2014 3782 2026 3834
rect 2078 3782 2090 3834
rect 2142 3782 2154 3834
rect 2206 3782 2218 3834
rect 2270 3782 3986 3834
rect 4038 3782 4050 3834
rect 4102 3782 4114 3834
rect 4166 3782 4178 3834
rect 4230 3782 4242 3834
rect 4294 3782 6010 3834
rect 6062 3782 6074 3834
rect 6126 3782 6138 3834
rect 6190 3782 6202 3834
rect 6254 3782 6266 3834
rect 6318 3782 8034 3834
rect 8086 3782 8098 3834
rect 8150 3782 8162 3834
rect 8214 3782 8226 3834
rect 8278 3782 8290 3834
rect 8342 3782 9200 3834
rect 1104 3760 9200 3782
rect 2314 3680 2320 3732
rect 2372 3680 2378 3732
rect 4614 3720 4620 3732
rect 4172 3692 4620 3720
rect 1949 3519 2007 3525
rect 1949 3485 1961 3519
rect 1995 3516 2007 3519
rect 2332 3516 2360 3680
rect 4065 3519 4123 3525
rect 4065 3516 4077 3519
rect 1995 3488 2360 3516
rect 3988 3488 4077 3516
rect 1995 3485 2007 3488
rect 1949 3479 2007 3485
rect 3988 3460 4016 3488
rect 4065 3485 4077 3488
rect 4111 3485 4123 3519
rect 4172 3516 4200 3692
rect 4614 3680 4620 3692
rect 4672 3720 4678 3732
rect 4672 3692 5120 3720
rect 4672 3680 4678 3692
rect 4246 3612 4252 3664
rect 4304 3652 4310 3664
rect 4801 3655 4859 3661
rect 4801 3652 4813 3655
rect 4304 3624 4813 3652
rect 4304 3612 4310 3624
rect 4801 3621 4813 3624
rect 4847 3621 4859 3655
rect 4801 3615 4859 3621
rect 4341 3587 4399 3593
rect 4341 3553 4353 3587
rect 4387 3584 4399 3587
rect 4525 3587 4583 3593
rect 4525 3584 4537 3587
rect 4387 3556 4537 3584
rect 4387 3553 4399 3556
rect 4341 3547 4399 3553
rect 4525 3553 4537 3556
rect 4571 3584 4583 3587
rect 4706 3584 4712 3596
rect 4571 3556 4712 3584
rect 4571 3553 4583 3556
rect 4525 3547 4583 3553
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 5092 3584 5120 3692
rect 5166 3680 5172 3732
rect 5224 3680 5230 3732
rect 7742 3680 7748 3732
rect 7800 3680 7806 3732
rect 5442 3584 5448 3596
rect 5092 3556 5448 3584
rect 5442 3544 5448 3556
rect 5500 3584 5506 3596
rect 5721 3587 5779 3593
rect 5721 3584 5733 3587
rect 5500 3556 5733 3584
rect 5500 3544 5506 3556
rect 5721 3553 5733 3556
rect 5767 3553 5779 3587
rect 7760 3584 7788 3680
rect 8662 3612 8668 3664
rect 8720 3612 8726 3664
rect 7760 3556 8064 3584
rect 5721 3547 5779 3553
rect 4249 3519 4307 3525
rect 4249 3516 4261 3519
rect 4172 3488 4261 3516
rect 4065 3479 4123 3485
rect 4249 3485 4261 3488
rect 4295 3485 4307 3519
rect 4249 3479 4307 3485
rect 4433 3519 4491 3525
rect 4433 3485 4445 3519
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 3970 3408 3976 3460
rect 4028 3448 4034 3460
rect 4448 3448 4476 3479
rect 4028 3420 4476 3448
rect 4724 3448 4752 3544
rect 5905 3519 5963 3525
rect 5905 3485 5917 3519
rect 5951 3516 5963 3519
rect 5951 3488 6408 3516
rect 5951 3485 5963 3488
rect 5905 3479 5963 3485
rect 6380 3460 6408 3488
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8036 3525 8064 3556
rect 7837 3519 7895 3525
rect 7837 3516 7849 3519
rect 7708 3488 7849 3516
rect 7708 3476 7714 3488
rect 7837 3485 7849 3488
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 8021 3519 8079 3525
rect 8021 3485 8033 3519
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 8202 3476 8208 3528
rect 8260 3516 8266 3528
rect 8481 3519 8539 3525
rect 8481 3516 8493 3519
rect 8260 3488 8493 3516
rect 8260 3476 8266 3488
rect 8481 3485 8493 3488
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 6150 3451 6208 3457
rect 6150 3448 6162 3451
rect 4724 3420 6162 3448
rect 4028 3408 4034 3420
rect 1670 3340 1676 3392
rect 1728 3380 1734 3392
rect 1765 3383 1823 3389
rect 1765 3380 1777 3383
rect 1728 3352 1777 3380
rect 1728 3340 1734 3352
rect 1765 3349 1777 3352
rect 1811 3349 1823 3383
rect 1765 3343 1823 3349
rect 3881 3383 3939 3389
rect 3881 3349 3893 3383
rect 3927 3380 3939 3383
rect 4338 3380 4344 3392
rect 3927 3352 4344 3380
rect 3927 3349 3939 3352
rect 3881 3343 3939 3349
rect 4338 3340 4344 3352
rect 4396 3340 4402 3392
rect 4448 3380 4476 3420
rect 6150 3417 6162 3420
rect 6196 3417 6208 3451
rect 6150 3411 6208 3417
rect 6362 3408 6368 3460
rect 6420 3408 6426 3460
rect 4890 3380 4896 3392
rect 4448 3352 4896 3380
rect 4890 3340 4896 3352
rect 4948 3340 4954 3392
rect 7285 3383 7343 3389
rect 7285 3349 7297 3383
rect 7331 3380 7343 3383
rect 7668 3380 7696 3476
rect 7331 3352 7696 3380
rect 7331 3349 7343 3352
rect 7285 3343 7343 3349
rect 7834 3340 7840 3392
rect 7892 3380 7898 3392
rect 7929 3383 7987 3389
rect 7929 3380 7941 3383
rect 7892 3352 7941 3380
rect 7892 3340 7898 3352
rect 7929 3349 7941 3352
rect 7975 3349 7987 3383
rect 7929 3343 7987 3349
rect 1104 3290 9200 3312
rect 1104 3238 2622 3290
rect 2674 3238 2686 3290
rect 2738 3238 2750 3290
rect 2802 3238 2814 3290
rect 2866 3238 2878 3290
rect 2930 3238 4646 3290
rect 4698 3238 4710 3290
rect 4762 3238 4774 3290
rect 4826 3238 4838 3290
rect 4890 3238 4902 3290
rect 4954 3238 6670 3290
rect 6722 3238 6734 3290
rect 6786 3238 6798 3290
rect 6850 3238 6862 3290
rect 6914 3238 6926 3290
rect 6978 3238 8694 3290
rect 8746 3238 8758 3290
rect 8810 3238 8822 3290
rect 8874 3238 8886 3290
rect 8938 3238 8950 3290
rect 9002 3238 9200 3290
rect 1104 3216 9200 3238
rect 2777 3179 2835 3185
rect 2777 3145 2789 3179
rect 2823 3176 2835 3179
rect 3142 3176 3148 3188
rect 2823 3148 3148 3176
rect 2823 3145 2835 3148
rect 2777 3139 2835 3145
rect 3142 3136 3148 3148
rect 3200 3136 3206 3188
rect 5442 3136 5448 3188
rect 5500 3176 5506 3188
rect 6089 3179 6147 3185
rect 6089 3176 6101 3179
rect 5500 3148 6101 3176
rect 5500 3136 5506 3148
rect 6089 3145 6101 3148
rect 6135 3145 6147 3179
rect 6089 3139 6147 3145
rect 2590 3108 2596 3120
rect 1412 3080 2596 3108
rect 1412 3052 1440 3080
rect 2590 3068 2596 3080
rect 2648 3108 2654 3120
rect 4617 3111 4675 3117
rect 2648 3080 2774 3108
rect 2648 3068 2654 3080
rect 1394 3000 1400 3052
rect 1452 3000 1458 3052
rect 1670 3049 1676 3052
rect 1664 3040 1676 3049
rect 1631 3012 1676 3040
rect 1664 3003 1676 3012
rect 1670 3000 1676 3003
rect 1728 3000 1734 3052
rect 2746 2972 2774 3080
rect 4617 3077 4629 3111
rect 4663 3108 4675 3111
rect 5074 3108 5080 3120
rect 4663 3080 5080 3108
rect 4663 3077 4675 3080
rect 4617 3071 4675 3077
rect 5074 3068 5080 3080
rect 5132 3068 5138 3120
rect 6104 3108 6132 3139
rect 7742 3136 7748 3188
rect 7800 3136 7806 3188
rect 6610 3111 6668 3117
rect 6610 3108 6622 3111
rect 6104 3080 6622 3108
rect 6610 3077 6622 3080
rect 6656 3077 6668 3111
rect 6610 3071 6668 3077
rect 4430 3000 4436 3052
rect 4488 3000 4494 3052
rect 4982 3049 4988 3052
rect 4976 3040 4988 3049
rect 4943 3012 4988 3040
rect 4976 3003 4988 3012
rect 4982 3000 4988 3003
rect 5040 3000 5046 3052
rect 6362 3000 6368 3052
rect 6420 3000 6426 3052
rect 7760 3040 7788 3136
rect 7834 3068 7840 3120
rect 7892 3108 7898 3120
rect 8205 3111 8263 3117
rect 7892 3080 8156 3108
rect 7892 3068 7898 3080
rect 8021 3043 8079 3049
rect 8021 3040 8033 3043
rect 7760 3012 8033 3040
rect 8021 3009 8033 3012
rect 8067 3009 8079 3043
rect 8128 3040 8156 3080
rect 8205 3077 8217 3111
rect 8251 3108 8263 3111
rect 8481 3111 8539 3117
rect 8481 3108 8493 3111
rect 8251 3080 8493 3108
rect 8251 3077 8263 3080
rect 8205 3071 8263 3077
rect 8481 3077 8493 3080
rect 8527 3077 8539 3111
rect 8481 3071 8539 3077
rect 8297 3043 8355 3049
rect 8297 3040 8309 3043
rect 8128 3012 8309 3040
rect 8021 3003 8079 3009
rect 8297 3009 8309 3012
rect 8343 3009 8355 3043
rect 8297 3003 8355 3009
rect 4448 2972 4476 3000
rect 4709 2975 4767 2981
rect 4709 2972 4721 2975
rect 2746 2944 4721 2972
rect 3344 2913 3372 2944
rect 4709 2941 4721 2944
rect 4755 2941 4767 2975
rect 4709 2935 4767 2941
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 7837 2975 7895 2981
rect 7837 2972 7849 2975
rect 7800 2944 7849 2972
rect 7800 2932 7806 2944
rect 7837 2941 7849 2944
rect 7883 2941 7895 2975
rect 7837 2935 7895 2941
rect 3329 2907 3387 2913
rect 3329 2873 3341 2907
rect 3375 2873 3387 2907
rect 3329 2867 3387 2873
rect 4246 2864 4252 2916
rect 4304 2904 4310 2916
rect 4430 2904 4436 2916
rect 4304 2876 4436 2904
rect 4304 2864 4310 2876
rect 4430 2864 4436 2876
rect 4488 2864 4494 2916
rect 7834 2796 7840 2848
rect 7892 2836 7898 2848
rect 8665 2839 8723 2845
rect 8665 2836 8677 2839
rect 7892 2808 8677 2836
rect 7892 2796 7898 2808
rect 8665 2805 8677 2808
rect 8711 2805 8723 2839
rect 8665 2799 8723 2805
rect 1104 2746 9200 2768
rect 1104 2694 1962 2746
rect 2014 2694 2026 2746
rect 2078 2694 2090 2746
rect 2142 2694 2154 2746
rect 2206 2694 2218 2746
rect 2270 2694 3986 2746
rect 4038 2694 4050 2746
rect 4102 2694 4114 2746
rect 4166 2694 4178 2746
rect 4230 2694 4242 2746
rect 4294 2694 6010 2746
rect 6062 2694 6074 2746
rect 6126 2694 6138 2746
rect 6190 2694 6202 2746
rect 6254 2694 6266 2746
rect 6318 2694 8034 2746
rect 8086 2694 8098 2746
rect 8150 2694 8162 2746
rect 8214 2694 8226 2746
rect 8278 2694 8290 2746
rect 8342 2694 9200 2746
rect 1104 2672 9200 2694
rect 2590 2632 2596 2644
rect 2240 2604 2596 2632
rect 2240 2505 2268 2604
rect 2590 2592 2596 2604
rect 2648 2592 2654 2644
rect 3605 2635 3663 2641
rect 3605 2601 3617 2635
rect 3651 2632 3663 2635
rect 3786 2632 3792 2644
rect 3651 2604 3792 2632
rect 3651 2601 3663 2604
rect 3605 2595 3663 2601
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 4338 2592 4344 2644
rect 4396 2592 4402 2644
rect 4522 2592 4528 2644
rect 4580 2632 4586 2644
rect 4617 2635 4675 2641
rect 4617 2632 4629 2635
rect 4580 2604 4629 2632
rect 4580 2592 4586 2604
rect 4617 2601 4629 2604
rect 4663 2601 4675 2635
rect 4617 2595 4675 2601
rect 7926 2592 7932 2644
rect 7984 2632 7990 2644
rect 8021 2635 8079 2641
rect 8021 2632 8033 2635
rect 7984 2604 8033 2632
rect 7984 2592 7990 2604
rect 8021 2601 8033 2604
rect 8067 2601 8079 2635
rect 8021 2595 8079 2601
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 8754 2632 8760 2644
rect 8711 2604 8760 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 8754 2592 8760 2604
rect 8812 2592 8818 2644
rect 3881 2567 3939 2573
rect 3881 2533 3893 2567
rect 3927 2533 3939 2567
rect 3881 2527 3939 2533
rect 2225 2499 2283 2505
rect 2225 2465 2237 2499
rect 2271 2465 2283 2499
rect 2225 2459 2283 2465
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2428 2007 2431
rect 3896 2428 3924 2527
rect 7742 2456 7748 2508
rect 7800 2496 7806 2508
rect 7800 2468 7972 2496
rect 7800 2456 7806 2468
rect 1995 2400 3924 2428
rect 4157 2431 4215 2437
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 4157 2397 4169 2431
rect 4203 2397 4215 2431
rect 4157 2391 4215 2397
rect 2470 2363 2528 2369
rect 2470 2360 2482 2363
rect 2148 2332 2482 2360
rect 2148 2301 2176 2332
rect 2470 2329 2482 2332
rect 2516 2329 2528 2363
rect 2470 2323 2528 2329
rect 2590 2320 2596 2372
rect 2648 2360 2654 2372
rect 4172 2360 4200 2391
rect 4430 2388 4436 2440
rect 4488 2388 4494 2440
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2428 4951 2431
rect 5166 2428 5172 2440
rect 4939 2400 5172 2428
rect 4939 2397 4951 2400
rect 4893 2391 4951 2397
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5350 2388 5356 2440
rect 5408 2388 5414 2440
rect 7653 2431 7711 2437
rect 7653 2397 7665 2431
rect 7699 2428 7711 2431
rect 7834 2428 7840 2440
rect 7699 2400 7840 2428
rect 7699 2397 7711 2400
rect 7653 2391 7711 2397
rect 7834 2388 7840 2400
rect 7892 2388 7898 2440
rect 7944 2437 7972 2468
rect 7929 2431 7987 2437
rect 7929 2397 7941 2431
rect 7975 2397 7987 2431
rect 7929 2391 7987 2397
rect 4617 2363 4675 2369
rect 4617 2360 4629 2363
rect 2648 2332 4629 2360
rect 2648 2320 2654 2332
rect 4617 2329 4629 2332
rect 4663 2329 4675 2363
rect 4617 2323 4675 2329
rect 4801 2363 4859 2369
rect 4801 2329 4813 2363
rect 4847 2360 4859 2363
rect 5368 2360 5396 2388
rect 8389 2363 8447 2369
rect 8389 2360 8401 2363
rect 4847 2332 5396 2360
rect 7852 2332 8401 2360
rect 4847 2329 4859 2332
rect 4801 2323 4859 2329
rect 7852 2301 7880 2332
rect 8389 2329 8401 2332
rect 8435 2329 8447 2363
rect 8389 2323 8447 2329
rect 2133 2295 2191 2301
rect 2133 2261 2145 2295
rect 2179 2261 2191 2295
rect 2133 2255 2191 2261
rect 7837 2295 7895 2301
rect 7837 2261 7849 2295
rect 7883 2261 7895 2295
rect 7837 2255 7895 2261
rect 1104 2202 9200 2224
rect 1104 2150 2622 2202
rect 2674 2150 2686 2202
rect 2738 2150 2750 2202
rect 2802 2150 2814 2202
rect 2866 2150 2878 2202
rect 2930 2150 4646 2202
rect 4698 2150 4710 2202
rect 4762 2150 4774 2202
rect 4826 2150 4838 2202
rect 4890 2150 4902 2202
rect 4954 2150 6670 2202
rect 6722 2150 6734 2202
rect 6786 2150 6798 2202
rect 6850 2150 6862 2202
rect 6914 2150 6926 2202
rect 6978 2150 8694 2202
rect 8746 2150 8758 2202
rect 8810 2150 8822 2202
rect 8874 2150 8886 2202
rect 8938 2150 8950 2202
rect 9002 2150 9200 2202
rect 1104 2128 9200 2150
<< via1 >>
rect 2622 9766 2674 9818
rect 2686 9766 2738 9818
rect 2750 9766 2802 9818
rect 2814 9766 2866 9818
rect 2878 9766 2930 9818
rect 4646 9766 4698 9818
rect 4710 9766 4762 9818
rect 4774 9766 4826 9818
rect 4838 9766 4890 9818
rect 4902 9766 4954 9818
rect 6670 9766 6722 9818
rect 6734 9766 6786 9818
rect 6798 9766 6850 9818
rect 6862 9766 6914 9818
rect 6926 9766 6978 9818
rect 8694 9766 8746 9818
rect 8758 9766 8810 9818
rect 8822 9766 8874 9818
rect 8886 9766 8938 9818
rect 8950 9766 9002 9818
rect 5816 9596 5868 9648
rect 6368 9435 6420 9444
rect 6368 9401 6377 9435
rect 6377 9401 6411 9435
rect 6411 9401 6420 9435
rect 6368 9392 6420 9401
rect 1962 9222 2014 9274
rect 2026 9222 2078 9274
rect 2090 9222 2142 9274
rect 2154 9222 2206 9274
rect 2218 9222 2270 9274
rect 3986 9222 4038 9274
rect 4050 9222 4102 9274
rect 4114 9222 4166 9274
rect 4178 9222 4230 9274
rect 4242 9222 4294 9274
rect 6010 9222 6062 9274
rect 6074 9222 6126 9274
rect 6138 9222 6190 9274
rect 6202 9222 6254 9274
rect 6266 9222 6318 9274
rect 8034 9222 8086 9274
rect 8098 9222 8150 9274
rect 8162 9222 8214 9274
rect 8226 9222 8278 9274
rect 8290 9222 8342 9274
rect 6368 9120 6420 9172
rect 1492 8916 1544 8968
rect 2964 8848 3016 8900
rect 4344 8959 4396 8968
rect 4344 8925 4353 8959
rect 4353 8925 4387 8959
rect 4387 8925 4396 8959
rect 4344 8916 4396 8925
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 8668 9095 8720 9104
rect 8668 9061 8677 9095
rect 8677 9061 8711 9095
rect 8711 9061 8720 9095
rect 8668 9052 8720 9061
rect 7748 9027 7800 9036
rect 7748 8993 7757 9027
rect 7757 8993 7791 9027
rect 7791 8993 7800 9027
rect 7748 8984 7800 8993
rect 5724 8848 5776 8900
rect 5816 8848 5868 8900
rect 3056 8780 3108 8832
rect 3424 8780 3476 8832
rect 5632 8780 5684 8832
rect 2622 8678 2674 8730
rect 2686 8678 2738 8730
rect 2750 8678 2802 8730
rect 2814 8678 2866 8730
rect 2878 8678 2930 8730
rect 4646 8678 4698 8730
rect 4710 8678 4762 8730
rect 4774 8678 4826 8730
rect 4838 8678 4890 8730
rect 4902 8678 4954 8730
rect 6670 8678 6722 8730
rect 6734 8678 6786 8730
rect 6798 8678 6850 8730
rect 6862 8678 6914 8730
rect 6926 8678 6978 8730
rect 8694 8678 8746 8730
rect 8758 8678 8810 8730
rect 8822 8678 8874 8730
rect 8886 8678 8938 8730
rect 8950 8678 9002 8730
rect 2964 8619 3016 8628
rect 2964 8585 2973 8619
rect 2973 8585 3007 8619
rect 3007 8585 3016 8619
rect 2964 8576 3016 8585
rect 3424 8576 3476 8628
rect 5724 8619 5776 8628
rect 5724 8585 5733 8619
rect 5733 8585 5767 8619
rect 5767 8585 5776 8619
rect 5724 8576 5776 8585
rect 1492 8440 1544 8492
rect 1676 8483 1728 8492
rect 1676 8449 1710 8483
rect 1710 8449 1728 8483
rect 1676 8440 1728 8449
rect 2504 8440 2556 8492
rect 5080 8440 5132 8492
rect 5632 8440 5684 8492
rect 5724 8440 5776 8492
rect 6368 8483 6420 8492
rect 6368 8449 6377 8483
rect 6377 8449 6411 8483
rect 6411 8449 6420 8483
rect 6368 8440 6420 8449
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 3240 8236 3292 8288
rect 3424 8236 3476 8288
rect 4528 8236 4580 8288
rect 4620 8279 4672 8288
rect 4620 8245 4629 8279
rect 4629 8245 4663 8279
rect 4663 8245 4672 8279
rect 4620 8236 4672 8245
rect 4988 8279 5040 8288
rect 4988 8245 4997 8279
rect 4997 8245 5031 8279
rect 5031 8245 5040 8279
rect 4988 8236 5040 8245
rect 7932 8236 7984 8288
rect 1962 8134 2014 8186
rect 2026 8134 2078 8186
rect 2090 8134 2142 8186
rect 2154 8134 2206 8186
rect 2218 8134 2270 8186
rect 3986 8134 4038 8186
rect 4050 8134 4102 8186
rect 4114 8134 4166 8186
rect 4178 8134 4230 8186
rect 4242 8134 4294 8186
rect 6010 8134 6062 8186
rect 6074 8134 6126 8186
rect 6138 8134 6190 8186
rect 6202 8134 6254 8186
rect 6266 8134 6318 8186
rect 8034 8134 8086 8186
rect 8098 8134 8150 8186
rect 8162 8134 8214 8186
rect 8226 8134 8278 8186
rect 8290 8134 8342 8186
rect 1676 8032 1728 8084
rect 3516 7964 3568 8016
rect 4988 8032 5040 8084
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 1400 7871 1452 7880
rect 1400 7837 1409 7871
rect 1409 7837 1443 7871
rect 1443 7837 1452 7871
rect 1400 7828 1452 7837
rect 2228 7871 2280 7880
rect 2228 7837 2237 7871
rect 2237 7837 2271 7871
rect 2271 7837 2280 7871
rect 2228 7828 2280 7837
rect 3240 7871 3292 7880
rect 3240 7837 3249 7871
rect 3249 7837 3283 7871
rect 3283 7837 3292 7871
rect 3240 7828 3292 7837
rect 3424 7871 3476 7880
rect 3424 7837 3433 7871
rect 3433 7837 3467 7871
rect 3467 7837 3476 7871
rect 3424 7828 3476 7837
rect 3516 7828 3568 7880
rect 4620 7828 4672 7880
rect 3700 7760 3752 7812
rect 4160 7760 4212 7812
rect 4344 7760 4396 7812
rect 4436 7760 4488 7812
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 5816 7871 5868 7880
rect 5816 7837 5825 7871
rect 5825 7837 5859 7871
rect 5859 7837 5868 7871
rect 5816 7828 5868 7837
rect 5908 7828 5960 7880
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 9128 7692 9180 7744
rect 2622 7590 2674 7642
rect 2686 7590 2738 7642
rect 2750 7590 2802 7642
rect 2814 7590 2866 7642
rect 2878 7590 2930 7642
rect 4646 7590 4698 7642
rect 4710 7590 4762 7642
rect 4774 7590 4826 7642
rect 4838 7590 4890 7642
rect 4902 7590 4954 7642
rect 6670 7590 6722 7642
rect 6734 7590 6786 7642
rect 6798 7590 6850 7642
rect 6862 7590 6914 7642
rect 6926 7590 6978 7642
rect 8694 7590 8746 7642
rect 8758 7590 8810 7642
rect 8822 7590 8874 7642
rect 8886 7590 8938 7642
rect 8950 7590 9002 7642
rect 2228 7488 2280 7540
rect 2504 7488 2556 7540
rect 3240 7488 3292 7540
rect 5724 7488 5776 7540
rect 5816 7488 5868 7540
rect 7748 7488 7800 7540
rect 7932 7488 7984 7540
rect 3056 7352 3108 7404
rect 3240 7352 3292 7404
rect 3608 7284 3660 7336
rect 3884 7284 3936 7336
rect 4436 7420 4488 7472
rect 4528 7420 4580 7472
rect 4344 7395 4396 7404
rect 4344 7361 4353 7395
rect 4353 7361 4387 7395
rect 4387 7361 4396 7395
rect 4344 7352 4396 7361
rect 3424 7216 3476 7268
rect 3332 7148 3384 7200
rect 4068 7216 4120 7268
rect 5908 7352 5960 7404
rect 6000 7395 6052 7404
rect 6000 7361 6009 7395
rect 6009 7361 6043 7395
rect 6043 7361 6052 7395
rect 6000 7352 6052 7361
rect 6368 7395 6420 7404
rect 6368 7361 6377 7395
rect 6377 7361 6411 7395
rect 6411 7361 6420 7395
rect 6368 7352 6420 7361
rect 5632 7284 5684 7336
rect 7380 7352 7432 7404
rect 4344 7148 4396 7200
rect 5448 7148 5500 7200
rect 5632 7148 5684 7200
rect 8392 7259 8444 7268
rect 8392 7225 8401 7259
rect 8401 7225 8435 7259
rect 8435 7225 8444 7259
rect 8392 7216 8444 7225
rect 5816 7148 5868 7200
rect 6000 7148 6052 7200
rect 7748 7191 7800 7200
rect 7748 7157 7757 7191
rect 7757 7157 7791 7191
rect 7791 7157 7800 7191
rect 7748 7148 7800 7157
rect 1962 7046 2014 7098
rect 2026 7046 2078 7098
rect 2090 7046 2142 7098
rect 2154 7046 2206 7098
rect 2218 7046 2270 7098
rect 3986 7046 4038 7098
rect 4050 7046 4102 7098
rect 4114 7046 4166 7098
rect 4178 7046 4230 7098
rect 4242 7046 4294 7098
rect 6010 7046 6062 7098
rect 6074 7046 6126 7098
rect 6138 7046 6190 7098
rect 6202 7046 6254 7098
rect 6266 7046 6318 7098
rect 8034 7046 8086 7098
rect 8098 7046 8150 7098
rect 8162 7046 8214 7098
rect 8226 7046 8278 7098
rect 8290 7046 8342 7098
rect 3700 6944 3752 6996
rect 5448 6944 5500 6996
rect 8484 6944 8536 6996
rect 3332 6740 3384 6792
rect 3424 6783 3476 6792
rect 3424 6749 3433 6783
rect 3433 6749 3467 6783
rect 3467 6749 3476 6783
rect 3424 6740 3476 6749
rect 5356 6876 5408 6928
rect 3608 6783 3660 6792
rect 3608 6749 3617 6783
rect 3617 6749 3651 6783
rect 3651 6749 3660 6783
rect 3608 6740 3660 6749
rect 3700 6740 3752 6792
rect 3884 6740 3936 6792
rect 4068 6740 4120 6792
rect 4436 6808 4488 6860
rect 7472 6919 7524 6928
rect 7472 6885 7481 6919
rect 7481 6885 7515 6919
rect 7515 6885 7524 6919
rect 7472 6876 7524 6885
rect 4344 6783 4396 6792
rect 4344 6749 4353 6783
rect 4353 6749 4387 6783
rect 4387 6749 4396 6783
rect 4344 6740 4396 6749
rect 2504 6672 2556 6724
rect 6368 6740 6420 6792
rect 7932 6740 7984 6792
rect 8576 6808 8628 6860
rect 8484 6740 8536 6792
rect 5908 6672 5960 6724
rect 7380 6672 7432 6724
rect 7656 6672 7708 6724
rect 1492 6647 1544 6656
rect 1492 6613 1501 6647
rect 1501 6613 1535 6647
rect 1535 6613 1544 6647
rect 1492 6604 1544 6613
rect 3056 6604 3108 6656
rect 3700 6604 3752 6656
rect 3884 6647 3936 6656
rect 3884 6613 3893 6647
rect 3893 6613 3927 6647
rect 3927 6613 3936 6647
rect 3884 6604 3936 6613
rect 4068 6604 4120 6656
rect 4988 6604 5040 6656
rect 8392 6604 8444 6656
rect 2622 6502 2674 6554
rect 2686 6502 2738 6554
rect 2750 6502 2802 6554
rect 2814 6502 2866 6554
rect 2878 6502 2930 6554
rect 4646 6502 4698 6554
rect 4710 6502 4762 6554
rect 4774 6502 4826 6554
rect 4838 6502 4890 6554
rect 4902 6502 4954 6554
rect 6670 6502 6722 6554
rect 6734 6502 6786 6554
rect 6798 6502 6850 6554
rect 6862 6502 6914 6554
rect 6926 6502 6978 6554
rect 8694 6502 8746 6554
rect 8758 6502 8810 6554
rect 8822 6502 8874 6554
rect 8886 6502 8938 6554
rect 8950 6502 9002 6554
rect 1492 6400 1544 6452
rect 3332 6400 3384 6452
rect 3240 6264 3292 6316
rect 3608 6264 3660 6316
rect 5172 6400 5224 6452
rect 7472 6400 7524 6452
rect 4068 6332 4120 6384
rect 4344 6307 4396 6316
rect 4344 6273 4378 6307
rect 4378 6273 4396 6307
rect 4344 6264 4396 6273
rect 5816 6264 5868 6316
rect 8300 6332 8352 6384
rect 3148 6171 3200 6180
rect 3148 6137 3157 6171
rect 3157 6137 3191 6171
rect 3191 6137 3200 6171
rect 3148 6128 3200 6137
rect 3608 6128 3660 6180
rect 2412 6103 2464 6112
rect 2412 6069 2421 6103
rect 2421 6069 2455 6103
rect 2455 6069 2464 6103
rect 2412 6060 2464 6069
rect 2688 6103 2740 6112
rect 2688 6069 2697 6103
rect 2697 6069 2731 6103
rect 2731 6069 2740 6103
rect 2688 6060 2740 6069
rect 3056 6103 3108 6112
rect 3056 6069 3065 6103
rect 3065 6069 3099 6103
rect 3099 6069 3108 6103
rect 3056 6060 3108 6069
rect 3424 6060 3476 6112
rect 7380 6196 7432 6248
rect 4068 6060 4120 6112
rect 4436 6060 4488 6112
rect 8484 6196 8536 6248
rect 7840 6060 7892 6112
rect 7932 6103 7984 6112
rect 7932 6069 7941 6103
rect 7941 6069 7975 6103
rect 7975 6069 7984 6103
rect 7932 6060 7984 6069
rect 8024 6060 8076 6112
rect 1962 5958 2014 6010
rect 2026 5958 2078 6010
rect 2090 5958 2142 6010
rect 2154 5958 2206 6010
rect 2218 5958 2270 6010
rect 3986 5958 4038 6010
rect 4050 5958 4102 6010
rect 4114 5958 4166 6010
rect 4178 5958 4230 6010
rect 4242 5958 4294 6010
rect 6010 5958 6062 6010
rect 6074 5958 6126 6010
rect 6138 5958 6190 6010
rect 6202 5958 6254 6010
rect 6266 5958 6318 6010
rect 8034 5958 8086 6010
rect 8098 5958 8150 6010
rect 8162 5958 8214 6010
rect 8226 5958 8278 6010
rect 8290 5958 8342 6010
rect 756 5856 808 5908
rect 2504 5856 2556 5908
rect 2688 5856 2740 5908
rect 1492 5720 1544 5772
rect 2412 5720 2464 5772
rect 3148 5856 3200 5908
rect 3240 5856 3292 5908
rect 3884 5856 3936 5908
rect 5080 5899 5132 5908
rect 5080 5865 5089 5899
rect 5089 5865 5123 5899
rect 5123 5865 5132 5899
rect 5080 5856 5132 5865
rect 7932 5856 7984 5908
rect 8668 5899 8720 5908
rect 8668 5865 8677 5899
rect 8677 5865 8711 5899
rect 8711 5865 8720 5899
rect 8668 5856 8720 5865
rect 3424 5720 3476 5772
rect 3056 5652 3108 5704
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 7656 5695 7708 5704
rect 7656 5661 7665 5695
rect 7665 5661 7699 5695
rect 7699 5661 7708 5695
rect 7656 5652 7708 5661
rect 3700 5584 3752 5636
rect 7932 5584 7984 5636
rect 2412 5516 2464 5568
rect 5632 5559 5684 5568
rect 5632 5525 5641 5559
rect 5641 5525 5675 5559
rect 5675 5525 5684 5559
rect 5632 5516 5684 5525
rect 8300 5516 8352 5568
rect 2622 5414 2674 5466
rect 2686 5414 2738 5466
rect 2750 5414 2802 5466
rect 2814 5414 2866 5466
rect 2878 5414 2930 5466
rect 4646 5414 4698 5466
rect 4710 5414 4762 5466
rect 4774 5414 4826 5466
rect 4838 5414 4890 5466
rect 4902 5414 4954 5466
rect 6670 5414 6722 5466
rect 6734 5414 6786 5466
rect 6798 5414 6850 5466
rect 6862 5414 6914 5466
rect 6926 5414 6978 5466
rect 8694 5414 8746 5466
rect 8758 5414 8810 5466
rect 8822 5414 8874 5466
rect 8886 5414 8938 5466
rect 8950 5414 9002 5466
rect 3700 5355 3752 5364
rect 3700 5321 3709 5355
rect 3709 5321 3743 5355
rect 3743 5321 3752 5355
rect 3700 5312 3752 5321
rect 4344 5312 4396 5364
rect 5172 5312 5224 5364
rect 3056 5244 3108 5296
rect 2412 5219 2464 5228
rect 2412 5185 2421 5219
rect 2421 5185 2455 5219
rect 2455 5185 2464 5219
rect 2412 5176 2464 5185
rect 2504 5219 2556 5228
rect 2504 5185 2513 5219
rect 2513 5185 2547 5219
rect 2547 5185 2556 5219
rect 2504 5176 2556 5185
rect 3516 5219 3568 5228
rect 3516 5185 3525 5219
rect 3525 5185 3559 5219
rect 3559 5185 3568 5219
rect 3516 5176 3568 5185
rect 3884 5176 3936 5228
rect 5172 5176 5224 5228
rect 4436 5151 4488 5160
rect 4436 5117 4445 5151
rect 4445 5117 4479 5151
rect 4479 5117 4488 5151
rect 4436 5108 4488 5117
rect 1676 4972 1728 5024
rect 2780 4972 2832 5024
rect 4712 4972 4764 5024
rect 6184 5176 6236 5228
rect 7472 5176 7524 5228
rect 8300 5176 8352 5228
rect 6368 5151 6420 5160
rect 6368 5117 6377 5151
rect 6377 5117 6411 5151
rect 6411 5117 6420 5151
rect 6368 5108 6420 5117
rect 7840 5108 7892 5160
rect 7748 5015 7800 5024
rect 7748 4981 7757 5015
rect 7757 4981 7791 5015
rect 7791 4981 7800 5015
rect 7748 4972 7800 4981
rect 8392 4972 8444 5024
rect 8760 5015 8812 5024
rect 8760 4981 8769 5015
rect 8769 4981 8803 5015
rect 8803 4981 8812 5015
rect 8760 4972 8812 4981
rect 1962 4870 2014 4922
rect 2026 4870 2078 4922
rect 2090 4870 2142 4922
rect 2154 4870 2206 4922
rect 2218 4870 2270 4922
rect 3986 4870 4038 4922
rect 4050 4870 4102 4922
rect 4114 4870 4166 4922
rect 4178 4870 4230 4922
rect 4242 4870 4294 4922
rect 6010 4870 6062 4922
rect 6074 4870 6126 4922
rect 6138 4870 6190 4922
rect 6202 4870 6254 4922
rect 6266 4870 6318 4922
rect 8034 4870 8086 4922
rect 8098 4870 8150 4922
rect 8162 4870 8214 4922
rect 8226 4870 8278 4922
rect 8290 4870 8342 4922
rect 2780 4811 2832 4820
rect 2780 4777 2789 4811
rect 2789 4777 2823 4811
rect 2823 4777 2832 4811
rect 2780 4768 2832 4777
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 1676 4607 1728 4616
rect 1676 4573 1710 4607
rect 1710 4573 1728 4607
rect 1676 4564 1728 4573
rect 3148 4768 3200 4820
rect 3608 4768 3660 4820
rect 4528 4811 4580 4820
rect 4528 4777 4537 4811
rect 4537 4777 4571 4811
rect 4571 4777 4580 4811
rect 4528 4768 4580 4777
rect 5172 4768 5224 4820
rect 7656 4768 7708 4820
rect 8392 4768 8444 4820
rect 3056 4700 3108 4752
rect 3148 4564 3200 4616
rect 3424 4564 3476 4616
rect 3976 4607 4028 4616
rect 3976 4573 3985 4607
rect 3985 4573 4019 4607
rect 4019 4573 4028 4607
rect 3976 4564 4028 4573
rect 4344 4564 4396 4616
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 4896 4564 4948 4616
rect 6368 4564 6420 4616
rect 7472 4700 7524 4752
rect 7748 4607 7800 4616
rect 7748 4573 7757 4607
rect 7757 4573 7791 4607
rect 7791 4573 7800 4607
rect 7748 4564 7800 4573
rect 7840 4564 7892 4616
rect 4988 4496 5040 4548
rect 2964 4428 3016 4480
rect 3148 4428 3200 4480
rect 3516 4428 3568 4480
rect 3976 4428 4028 4480
rect 4344 4428 4396 4480
rect 5632 4428 5684 4480
rect 9128 4428 9180 4480
rect 2622 4326 2674 4378
rect 2686 4326 2738 4378
rect 2750 4326 2802 4378
rect 2814 4326 2866 4378
rect 2878 4326 2930 4378
rect 4646 4326 4698 4378
rect 4710 4326 4762 4378
rect 4774 4326 4826 4378
rect 4838 4326 4890 4378
rect 4902 4326 4954 4378
rect 6670 4326 6722 4378
rect 6734 4326 6786 4378
rect 6798 4326 6850 4378
rect 6862 4326 6914 4378
rect 6926 4326 6978 4378
rect 8694 4326 8746 4378
rect 8758 4326 8810 4378
rect 8822 4326 8874 4378
rect 8886 4326 8938 4378
rect 8950 4326 9002 4378
rect 3056 4224 3108 4276
rect 4252 4224 4304 4276
rect 4712 4224 4764 4276
rect 5172 4224 5224 4276
rect 7748 4224 7800 4276
rect 7564 4088 7616 4140
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 2504 4063 2556 4072
rect 2504 4029 2513 4063
rect 2513 4029 2547 4063
rect 2547 4029 2556 4063
rect 2504 4020 2556 4029
rect 4528 4020 4580 4072
rect 7932 4020 7984 4072
rect 2320 3884 2372 3936
rect 2964 3884 3016 3936
rect 4988 3927 5040 3936
rect 4988 3893 4997 3927
rect 4997 3893 5031 3927
rect 5031 3893 5040 3927
rect 4988 3884 5040 3893
rect 5172 3884 5224 3936
rect 7656 3884 7708 3936
rect 1962 3782 2014 3834
rect 2026 3782 2078 3834
rect 2090 3782 2142 3834
rect 2154 3782 2206 3834
rect 2218 3782 2270 3834
rect 3986 3782 4038 3834
rect 4050 3782 4102 3834
rect 4114 3782 4166 3834
rect 4178 3782 4230 3834
rect 4242 3782 4294 3834
rect 6010 3782 6062 3834
rect 6074 3782 6126 3834
rect 6138 3782 6190 3834
rect 6202 3782 6254 3834
rect 6266 3782 6318 3834
rect 8034 3782 8086 3834
rect 8098 3782 8150 3834
rect 8162 3782 8214 3834
rect 8226 3782 8278 3834
rect 8290 3782 8342 3834
rect 2320 3680 2372 3732
rect 4620 3723 4672 3732
rect 4620 3689 4629 3723
rect 4629 3689 4663 3723
rect 4663 3689 4672 3723
rect 4620 3680 4672 3689
rect 4252 3612 4304 3664
rect 4712 3544 4764 3596
rect 5172 3723 5224 3732
rect 5172 3689 5181 3723
rect 5181 3689 5215 3723
rect 5215 3689 5224 3723
rect 5172 3680 5224 3689
rect 7748 3680 7800 3732
rect 5448 3544 5500 3596
rect 8668 3655 8720 3664
rect 8668 3621 8677 3655
rect 8677 3621 8711 3655
rect 8711 3621 8720 3655
rect 8668 3612 8720 3621
rect 3976 3408 4028 3460
rect 7656 3476 7708 3528
rect 8208 3476 8260 3528
rect 1676 3340 1728 3392
rect 4344 3340 4396 3392
rect 6368 3408 6420 3460
rect 4896 3340 4948 3392
rect 7840 3340 7892 3392
rect 2622 3238 2674 3290
rect 2686 3238 2738 3290
rect 2750 3238 2802 3290
rect 2814 3238 2866 3290
rect 2878 3238 2930 3290
rect 4646 3238 4698 3290
rect 4710 3238 4762 3290
rect 4774 3238 4826 3290
rect 4838 3238 4890 3290
rect 4902 3238 4954 3290
rect 6670 3238 6722 3290
rect 6734 3238 6786 3290
rect 6798 3238 6850 3290
rect 6862 3238 6914 3290
rect 6926 3238 6978 3290
rect 8694 3238 8746 3290
rect 8758 3238 8810 3290
rect 8822 3238 8874 3290
rect 8886 3238 8938 3290
rect 8950 3238 9002 3290
rect 3148 3136 3200 3188
rect 5448 3136 5500 3188
rect 2596 3068 2648 3120
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 1676 3043 1728 3052
rect 1676 3009 1710 3043
rect 1710 3009 1728 3043
rect 1676 3000 1728 3009
rect 5080 3068 5132 3120
rect 7748 3179 7800 3188
rect 7748 3145 7757 3179
rect 7757 3145 7791 3179
rect 7791 3145 7800 3179
rect 7748 3136 7800 3145
rect 4436 3000 4488 3052
rect 4988 3043 5040 3052
rect 4988 3009 5022 3043
rect 5022 3009 5040 3043
rect 4988 3000 5040 3009
rect 6368 3043 6420 3052
rect 6368 3009 6377 3043
rect 6377 3009 6411 3043
rect 6411 3009 6420 3043
rect 6368 3000 6420 3009
rect 7840 3068 7892 3120
rect 7748 2932 7800 2984
rect 4252 2864 4304 2916
rect 4436 2864 4488 2916
rect 7840 2796 7892 2848
rect 1962 2694 2014 2746
rect 2026 2694 2078 2746
rect 2090 2694 2142 2746
rect 2154 2694 2206 2746
rect 2218 2694 2270 2746
rect 3986 2694 4038 2746
rect 4050 2694 4102 2746
rect 4114 2694 4166 2746
rect 4178 2694 4230 2746
rect 4242 2694 4294 2746
rect 6010 2694 6062 2746
rect 6074 2694 6126 2746
rect 6138 2694 6190 2746
rect 6202 2694 6254 2746
rect 6266 2694 6318 2746
rect 8034 2694 8086 2746
rect 8098 2694 8150 2746
rect 8162 2694 8214 2746
rect 8226 2694 8278 2746
rect 8290 2694 8342 2746
rect 2596 2592 2648 2644
rect 3792 2592 3844 2644
rect 4344 2635 4396 2644
rect 4344 2601 4353 2635
rect 4353 2601 4387 2635
rect 4387 2601 4396 2635
rect 4344 2592 4396 2601
rect 4528 2592 4580 2644
rect 7932 2592 7984 2644
rect 8760 2592 8812 2644
rect 7748 2456 7800 2508
rect 2596 2320 2648 2372
rect 4436 2431 4488 2440
rect 4436 2397 4445 2431
rect 4445 2397 4479 2431
rect 4479 2397 4488 2431
rect 4436 2388 4488 2397
rect 5172 2388 5224 2440
rect 5356 2388 5408 2440
rect 7840 2388 7892 2440
rect 2622 2150 2674 2202
rect 2686 2150 2738 2202
rect 2750 2150 2802 2202
rect 2814 2150 2866 2202
rect 2878 2150 2930 2202
rect 4646 2150 4698 2202
rect 4710 2150 4762 2202
rect 4774 2150 4826 2202
rect 4838 2150 4890 2202
rect 4902 2150 4954 2202
rect 6670 2150 6722 2202
rect 6734 2150 6786 2202
rect 6798 2150 6850 2202
rect 6862 2150 6914 2202
rect 6926 2150 6978 2202
rect 8694 2150 8746 2202
rect 8758 2150 8810 2202
rect 8822 2150 8874 2202
rect 8886 2150 8938 2202
rect 8950 2150 9002 2202
<< metal2 >>
rect 5814 11661 5870 12461
rect 2622 9820 2930 9829
rect 2622 9818 2628 9820
rect 2684 9818 2708 9820
rect 2764 9818 2788 9820
rect 2844 9818 2868 9820
rect 2924 9818 2930 9820
rect 2684 9766 2686 9818
rect 2866 9766 2868 9818
rect 2622 9764 2628 9766
rect 2684 9764 2708 9766
rect 2764 9764 2788 9766
rect 2844 9764 2868 9766
rect 2924 9764 2930 9766
rect 2622 9755 2930 9764
rect 4646 9820 4954 9829
rect 4646 9818 4652 9820
rect 4708 9818 4732 9820
rect 4788 9818 4812 9820
rect 4868 9818 4892 9820
rect 4948 9818 4954 9820
rect 4708 9766 4710 9818
rect 4890 9766 4892 9818
rect 4646 9764 4652 9766
rect 4708 9764 4732 9766
rect 4788 9764 4812 9766
rect 4868 9764 4892 9766
rect 4948 9764 4954 9766
rect 4646 9755 4954 9764
rect 5828 9654 5856 11661
rect 6670 9820 6978 9829
rect 6670 9818 6676 9820
rect 6732 9818 6756 9820
rect 6812 9818 6836 9820
rect 6892 9818 6916 9820
rect 6972 9818 6978 9820
rect 6732 9766 6734 9818
rect 6914 9766 6916 9818
rect 6670 9764 6676 9766
rect 6732 9764 6756 9766
rect 6812 9764 6836 9766
rect 6892 9764 6916 9766
rect 6972 9764 6978 9766
rect 6670 9755 6978 9764
rect 8694 9820 9002 9829
rect 8694 9818 8700 9820
rect 8756 9818 8780 9820
rect 8836 9818 8860 9820
rect 8916 9818 8940 9820
rect 8996 9818 9002 9820
rect 8756 9766 8758 9818
rect 8938 9766 8940 9818
rect 8694 9764 8700 9766
rect 8756 9764 8780 9766
rect 8836 9764 8860 9766
rect 8916 9764 8940 9766
rect 8996 9764 9002 9766
rect 8694 9755 9002 9764
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 6368 9444 6420 9450
rect 6368 9386 6420 9392
rect 1962 9276 2270 9285
rect 1962 9274 1968 9276
rect 2024 9274 2048 9276
rect 2104 9274 2128 9276
rect 2184 9274 2208 9276
rect 2264 9274 2270 9276
rect 2024 9222 2026 9274
rect 2206 9222 2208 9274
rect 1962 9220 1968 9222
rect 2024 9220 2048 9222
rect 2104 9220 2128 9222
rect 2184 9220 2208 9222
rect 2264 9220 2270 9222
rect 1962 9211 2270 9220
rect 3986 9276 4294 9285
rect 3986 9274 3992 9276
rect 4048 9274 4072 9276
rect 4128 9274 4152 9276
rect 4208 9274 4232 9276
rect 4288 9274 4294 9276
rect 4048 9222 4050 9274
rect 4230 9222 4232 9274
rect 3986 9220 3992 9222
rect 4048 9220 4072 9222
rect 4128 9220 4152 9222
rect 4208 9220 4232 9222
rect 4288 9220 4294 9222
rect 3986 9211 4294 9220
rect 6010 9276 6318 9285
rect 6010 9274 6016 9276
rect 6072 9274 6096 9276
rect 6152 9274 6176 9276
rect 6232 9274 6256 9276
rect 6312 9274 6318 9276
rect 6072 9222 6074 9274
rect 6254 9222 6256 9274
rect 6010 9220 6016 9222
rect 6072 9220 6096 9222
rect 6152 9220 6176 9222
rect 6232 9220 6256 9222
rect 6312 9220 6318 9222
rect 6010 9211 6318 9220
rect 6380 9178 6408 9386
rect 8034 9276 8342 9285
rect 8034 9274 8040 9276
rect 8096 9274 8120 9276
rect 8176 9274 8200 9276
rect 8256 9274 8280 9276
rect 8336 9274 8342 9276
rect 8096 9222 8098 9274
rect 8278 9222 8280 9274
rect 8034 9220 8040 9222
rect 8096 9220 8120 9222
rect 8176 9220 8200 9222
rect 8256 9220 8280 9222
rect 8336 9220 8342 9222
rect 8034 9211 8342 9220
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 1492 8968 1544 8974
rect 4344 8968 4396 8974
rect 1492 8910 1544 8916
rect 3790 8936 3846 8945
rect 1504 8498 1532 8910
rect 2964 8900 3016 8906
rect 4344 8910 4396 8916
rect 4528 8968 4580 8974
rect 4528 8910 4580 8916
rect 3790 8871 3846 8880
rect 2964 8842 3016 8848
rect 2622 8732 2930 8741
rect 2622 8730 2628 8732
rect 2684 8730 2708 8732
rect 2764 8730 2788 8732
rect 2844 8730 2868 8732
rect 2924 8730 2930 8732
rect 2684 8678 2686 8730
rect 2866 8678 2868 8730
rect 2622 8676 2628 8678
rect 2684 8676 2708 8678
rect 2764 8676 2788 8678
rect 2844 8676 2868 8678
rect 2924 8676 2930 8678
rect 2622 8667 2930 8676
rect 2976 8634 3004 8842
rect 3056 8832 3108 8838
rect 3056 8774 3108 8780
rect 3424 8832 3476 8838
rect 3424 8774 3476 8780
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 1688 8090 1716 8434
rect 1962 8188 2270 8197
rect 1962 8186 1968 8188
rect 2024 8186 2048 8188
rect 2104 8186 2128 8188
rect 2184 8186 2208 8188
rect 2264 8186 2270 8188
rect 2024 8134 2026 8186
rect 2206 8134 2208 8186
rect 1962 8132 1968 8134
rect 2024 8132 2048 8134
rect 2104 8132 2128 8134
rect 2184 8132 2208 8134
rect 2264 8132 2270 8134
rect 1962 8123 2270 8132
rect 1676 8084 1728 8090
rect 1676 8026 1728 8032
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 2228 7880 2280 7886
rect 2228 7822 2280 7828
rect 1412 7585 1440 7822
rect 1398 7576 1454 7585
rect 2240 7546 2268 7822
rect 2516 7546 2544 8434
rect 2622 7644 2930 7653
rect 2622 7642 2628 7644
rect 2684 7642 2708 7644
rect 2764 7642 2788 7644
rect 2844 7642 2868 7644
rect 2924 7642 2930 7644
rect 2684 7590 2686 7642
rect 2866 7590 2868 7642
rect 2622 7588 2628 7590
rect 2684 7588 2708 7590
rect 2764 7588 2788 7590
rect 2844 7588 2868 7590
rect 2924 7588 2930 7590
rect 2622 7579 2930 7588
rect 1398 7511 1454 7520
rect 2228 7540 2280 7546
rect 2228 7482 2280 7488
rect 2504 7540 2556 7546
rect 2504 7482 2556 7488
rect 3068 7410 3096 8774
rect 3436 8634 3464 8774
rect 3424 8628 3476 8634
rect 3424 8570 3476 8576
rect 3240 8288 3292 8294
rect 3240 8230 3292 8236
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3252 7886 3280 8230
rect 3436 7886 3464 8230
rect 3516 8016 3568 8022
rect 3568 7964 3648 7970
rect 3516 7958 3648 7964
rect 3528 7942 3648 7958
rect 3240 7880 3292 7886
rect 3424 7880 3476 7886
rect 3240 7822 3292 7828
rect 3344 7828 3424 7834
rect 3516 7880 3568 7886
rect 3344 7822 3476 7828
rect 3514 7848 3516 7857
rect 3568 7848 3570 7857
rect 3252 7546 3280 7822
rect 3344 7806 3464 7822
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 3344 7426 3372 7806
rect 3514 7783 3570 7792
rect 3056 7404 3108 7410
rect 3056 7346 3108 7352
rect 3240 7404 3292 7410
rect 3344 7398 3464 7426
rect 3240 7346 3292 7352
rect 1962 7100 2270 7109
rect 1962 7098 1968 7100
rect 2024 7098 2048 7100
rect 2104 7098 2128 7100
rect 2184 7098 2208 7100
rect 2264 7098 2270 7100
rect 2024 7046 2026 7098
rect 2206 7046 2208 7098
rect 1962 7044 1968 7046
rect 2024 7044 2048 7046
rect 2104 7044 2128 7046
rect 2184 7044 2208 7046
rect 2264 7044 2270 7046
rect 1962 7035 2270 7044
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1504 6458 1532 6598
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 754 5944 810 5953
rect 754 5879 756 5888
rect 808 5879 810 5888
rect 756 5850 808 5856
rect 1504 5778 1532 6394
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 1962 6012 2270 6021
rect 1962 6010 1968 6012
rect 2024 6010 2048 6012
rect 2104 6010 2128 6012
rect 2184 6010 2208 6012
rect 2264 6010 2270 6012
rect 2024 5958 2026 6010
rect 2206 5958 2208 6010
rect 1962 5956 1968 5958
rect 2024 5956 2048 5958
rect 2104 5956 2128 5958
rect 2184 5956 2208 5958
rect 2264 5956 2270 5958
rect 1962 5947 2270 5956
rect 2424 5778 2452 6054
rect 2516 5914 2544 6666
rect 3056 6656 3108 6662
rect 3056 6598 3108 6604
rect 2622 6556 2930 6565
rect 2622 6554 2628 6556
rect 2684 6554 2708 6556
rect 2764 6554 2788 6556
rect 2844 6554 2868 6556
rect 2924 6554 2930 6556
rect 2684 6502 2686 6554
rect 2866 6502 2868 6554
rect 2622 6500 2628 6502
rect 2684 6500 2708 6502
rect 2764 6500 2788 6502
rect 2844 6500 2868 6502
rect 2924 6500 2930 6502
rect 2622 6491 2930 6500
rect 3068 6202 3096 6598
rect 3252 6322 3280 7346
rect 3436 7274 3464 7398
rect 3620 7342 3648 7942
rect 3700 7812 3752 7818
rect 3700 7754 3752 7760
rect 3608 7336 3660 7342
rect 3608 7278 3660 7284
rect 3424 7268 3476 7274
rect 3424 7210 3476 7216
rect 3332 7200 3384 7206
rect 3332 7142 3384 7148
rect 3344 6798 3372 7142
rect 3436 6798 3464 7210
rect 3712 7002 3740 7754
rect 3700 6996 3752 7002
rect 3700 6938 3752 6944
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3424 6792 3476 6798
rect 3424 6734 3476 6740
rect 3608 6792 3660 6798
rect 3608 6734 3660 6740
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3344 6458 3372 6734
rect 3332 6452 3384 6458
rect 3332 6394 3384 6400
rect 3240 6316 3292 6322
rect 3240 6258 3292 6264
rect 2976 6174 3096 6202
rect 3148 6180 3200 6186
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 2700 5914 2728 6054
rect 2504 5908 2556 5914
rect 2504 5850 2556 5856
rect 2688 5908 2740 5914
rect 2688 5850 2740 5856
rect 2976 5794 3004 6174
rect 3148 6122 3200 6128
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 1492 5772 1544 5778
rect 1492 5714 1544 5720
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2516 5766 3004 5794
rect 2412 5568 2464 5574
rect 2412 5510 2464 5516
rect 2424 5234 2452 5510
rect 2516 5234 2544 5766
rect 3068 5710 3096 6054
rect 3160 5914 3188 6122
rect 3252 5914 3280 6258
rect 3436 6118 3464 6734
rect 3620 6322 3648 6734
rect 3712 6662 3740 6734
rect 3700 6656 3752 6662
rect 3700 6598 3752 6604
rect 3608 6316 3660 6322
rect 3608 6258 3660 6264
rect 3608 6180 3660 6186
rect 3608 6122 3660 6128
rect 3424 6112 3476 6118
rect 3424 6054 3476 6060
rect 3148 5908 3200 5914
rect 3148 5850 3200 5856
rect 3240 5908 3292 5914
rect 3240 5850 3292 5856
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2622 5468 2930 5477
rect 2622 5466 2628 5468
rect 2684 5466 2708 5468
rect 2764 5466 2788 5468
rect 2844 5466 2868 5468
rect 2924 5466 2930 5468
rect 2684 5414 2686 5466
rect 2866 5414 2868 5466
rect 2622 5412 2628 5414
rect 2684 5412 2708 5414
rect 2764 5412 2788 5414
rect 2844 5412 2868 5414
rect 2924 5412 2930 5414
rect 2622 5403 2930 5412
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 2504 5228 2556 5234
rect 2504 5170 2556 5176
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1688 4622 1716 4966
rect 1962 4924 2270 4933
rect 1962 4922 1968 4924
rect 2024 4922 2048 4924
rect 2104 4922 2128 4924
rect 2184 4922 2208 4924
rect 2264 4922 2270 4924
rect 2024 4870 2026 4922
rect 2206 4870 2208 4922
rect 1962 4868 1968 4870
rect 2024 4868 2048 4870
rect 2104 4868 2128 4870
rect 2184 4868 2208 4870
rect 2264 4868 2270 4870
rect 1962 4859 2270 4868
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1412 3058 1440 4558
rect 2516 4078 2544 5170
rect 2780 5024 2832 5030
rect 2780 4966 2832 4972
rect 2792 4826 2820 4966
rect 2780 4820 2832 4826
rect 2780 4762 2832 4768
rect 3068 4758 3096 5238
rect 3160 4826 3188 5850
rect 3436 5778 3464 6054
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3056 4752 3108 4758
rect 3056 4694 3108 4700
rect 2964 4480 3016 4486
rect 2964 4422 3016 4428
rect 2622 4380 2930 4389
rect 2622 4378 2628 4380
rect 2684 4378 2708 4380
rect 2764 4378 2788 4380
rect 2844 4378 2868 4380
rect 2924 4378 2930 4380
rect 2684 4326 2686 4378
rect 2866 4326 2868 4378
rect 2622 4324 2628 4326
rect 2684 4324 2708 4326
rect 2764 4324 2788 4326
rect 2844 4324 2868 4326
rect 2924 4324 2930 4326
rect 2622 4315 2930 4324
rect 2504 4072 2556 4078
rect 2504 4014 2556 4020
rect 2320 3936 2372 3942
rect 2320 3878 2372 3884
rect 1962 3836 2270 3845
rect 1962 3834 1968 3836
rect 2024 3834 2048 3836
rect 2104 3834 2128 3836
rect 2184 3834 2208 3836
rect 2264 3834 2270 3836
rect 2024 3782 2026 3834
rect 2206 3782 2208 3834
rect 1962 3780 1968 3782
rect 2024 3780 2048 3782
rect 2104 3780 2128 3782
rect 2184 3780 2208 3782
rect 2264 3780 2270 3782
rect 1962 3771 2270 3780
rect 2332 3738 2360 3878
rect 2320 3732 2372 3738
rect 2320 3674 2372 3680
rect 1676 3392 1728 3398
rect 1676 3334 1728 3340
rect 1688 3058 1716 3334
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 1676 3052 1728 3058
rect 1676 2994 1728 3000
rect 1962 2748 2270 2757
rect 1962 2746 1968 2748
rect 2024 2746 2048 2748
rect 2104 2746 2128 2748
rect 2184 2746 2208 2748
rect 2264 2746 2270 2748
rect 2024 2694 2026 2746
rect 2206 2694 2208 2746
rect 1962 2692 1968 2694
rect 2024 2692 2048 2694
rect 2104 2692 2128 2694
rect 2184 2692 2208 2694
rect 2264 2692 2270 2694
rect 1962 2683 2270 2692
rect 2516 2530 2544 4014
rect 2976 3942 3004 4422
rect 3068 4282 3096 4694
rect 3436 4622 3464 5714
rect 3516 5228 3568 5234
rect 3516 5170 3568 5176
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3160 4486 3188 4558
rect 3528 4486 3556 5170
rect 3620 4826 3648 6122
rect 3804 5710 3832 8871
rect 3986 8188 4294 8197
rect 3986 8186 3992 8188
rect 4048 8186 4072 8188
rect 4128 8186 4152 8188
rect 4208 8186 4232 8188
rect 4288 8186 4294 8188
rect 4048 8134 4050 8186
rect 4230 8134 4232 8186
rect 3986 8132 3992 8134
rect 4048 8132 4072 8134
rect 4128 8132 4152 8134
rect 4208 8132 4232 8134
rect 4288 8132 4294 8134
rect 3986 8123 4294 8132
rect 4356 7818 4384 8910
rect 4540 8378 4568 8910
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 5632 8832 5684 8838
rect 5632 8774 5684 8780
rect 4646 8732 4954 8741
rect 4646 8730 4652 8732
rect 4708 8730 4732 8732
rect 4788 8730 4812 8732
rect 4868 8730 4892 8732
rect 4948 8730 4954 8732
rect 4708 8678 4710 8730
rect 4890 8678 4892 8730
rect 4646 8676 4652 8678
rect 4708 8676 4732 8678
rect 4788 8676 4812 8678
rect 4868 8676 4892 8678
rect 4948 8676 4954 8678
rect 4646 8667 4954 8676
rect 5644 8498 5672 8774
rect 5736 8634 5764 8842
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 5632 8492 5684 8498
rect 5632 8434 5684 8440
rect 5724 8492 5776 8498
rect 5724 8434 5776 8440
rect 4540 8350 4660 8378
rect 4632 8294 4660 8350
rect 4528 8288 4580 8294
rect 4528 8230 4580 8236
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 4434 7848 4490 7857
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 4344 7812 4396 7818
rect 4434 7783 4436 7792
rect 4344 7754 4396 7760
rect 4488 7783 4490 7792
rect 4436 7754 4488 7760
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 3896 6798 3924 7278
rect 4068 7268 4120 7274
rect 4172 7256 4200 7754
rect 4448 7562 4476 7754
rect 4356 7534 4476 7562
rect 4356 7410 4384 7534
rect 4540 7478 4568 8230
rect 4632 7886 4660 8230
rect 5000 8090 5028 8230
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4646 7644 4954 7653
rect 4646 7642 4652 7644
rect 4708 7642 4732 7644
rect 4788 7642 4812 7644
rect 4868 7642 4892 7644
rect 4948 7642 4954 7644
rect 4708 7590 4710 7642
rect 4890 7590 4892 7642
rect 4646 7588 4652 7590
rect 4708 7588 4732 7590
rect 4788 7588 4812 7590
rect 4868 7588 4892 7590
rect 4948 7588 4954 7590
rect 4646 7579 4954 7588
rect 4436 7472 4488 7478
rect 4436 7414 4488 7420
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4344 7404 4396 7410
rect 4344 7346 4396 7352
rect 4120 7228 4200 7256
rect 4068 7210 4120 7216
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 3986 7100 4294 7109
rect 3986 7098 3992 7100
rect 4048 7098 4072 7100
rect 4128 7098 4152 7100
rect 4208 7098 4232 7100
rect 4288 7098 4294 7100
rect 4048 7046 4050 7098
rect 4230 7046 4232 7098
rect 3986 7044 3992 7046
rect 4048 7044 4072 7046
rect 4128 7044 4152 7046
rect 4208 7044 4232 7046
rect 4288 7044 4294 7046
rect 3986 7035 4294 7044
rect 4356 6798 4384 7142
rect 4448 6866 4476 7414
rect 4436 6860 4488 6866
rect 4436 6802 4488 6808
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 4068 6792 4120 6798
rect 4068 6734 4120 6740
rect 4344 6792 4396 6798
rect 4344 6734 4396 6740
rect 4080 6662 4108 6734
rect 3884 6656 3936 6662
rect 3884 6598 3936 6604
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 3896 5914 3924 6598
rect 4646 6556 4954 6565
rect 4646 6554 4652 6556
rect 4708 6554 4732 6556
rect 4788 6554 4812 6556
rect 4868 6554 4892 6556
rect 4948 6554 4954 6556
rect 4708 6502 4710 6554
rect 4890 6502 4892 6554
rect 4646 6500 4652 6502
rect 4708 6500 4732 6502
rect 4788 6500 4812 6502
rect 4868 6500 4892 6502
rect 4948 6500 4954 6502
rect 4646 6491 4954 6500
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4080 6118 4108 6326
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3986 6012 4294 6021
rect 3986 6010 3992 6012
rect 4048 6010 4072 6012
rect 4128 6010 4152 6012
rect 4208 6010 4232 6012
rect 4288 6010 4294 6012
rect 4048 5958 4050 6010
rect 4230 5958 4232 6010
rect 3986 5956 3992 5958
rect 4048 5956 4072 5958
rect 4128 5956 4152 5958
rect 4208 5956 4232 5958
rect 4288 5956 4294 5958
rect 3986 5947 4294 5956
rect 3884 5908 3936 5914
rect 3884 5850 3936 5856
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3700 5636 3752 5642
rect 3700 5578 3752 5584
rect 3712 5370 3740 5578
rect 3700 5364 3752 5370
rect 3700 5306 3752 5312
rect 3896 5234 3924 5850
rect 4356 5370 4384 6258
rect 4436 6112 4488 6118
rect 4436 6054 4488 6060
rect 4344 5364 4396 5370
rect 4344 5306 4396 5312
rect 4448 5250 4476 6054
rect 4646 5468 4954 5477
rect 4646 5466 4652 5468
rect 4708 5466 4732 5468
rect 4788 5466 4812 5468
rect 4868 5466 4892 5468
rect 4948 5466 4954 5468
rect 4708 5414 4710 5466
rect 4890 5414 4892 5466
rect 4646 5412 4652 5414
rect 4708 5412 4732 5414
rect 4788 5412 4812 5414
rect 4868 5412 4892 5414
rect 4948 5412 4954 5414
rect 4646 5403 4954 5412
rect 5000 5250 5028 6598
rect 5092 5914 5120 8434
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5552 8090 5580 8366
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5368 6934 5396 7686
rect 5448 7200 5500 7206
rect 5448 7142 5500 7148
rect 5552 7154 5580 8026
rect 5644 7886 5672 8434
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5644 7342 5672 7822
rect 5736 7546 5764 8434
rect 5828 7886 5856 8842
rect 6380 8498 6408 9114
rect 8668 9104 8720 9110
rect 8668 9046 8720 9052
rect 7748 9036 7800 9042
rect 7748 8978 7800 8984
rect 6670 8732 6978 8741
rect 6670 8730 6676 8732
rect 6732 8730 6756 8732
rect 6812 8730 6836 8732
rect 6892 8730 6916 8732
rect 6972 8730 6978 8732
rect 6732 8678 6734 8730
rect 6914 8678 6916 8730
rect 6670 8676 6676 8678
rect 6732 8676 6756 8678
rect 6812 8676 6836 8678
rect 6892 8676 6916 8678
rect 6972 8676 6978 8678
rect 6670 8667 6978 8676
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6010 8188 6318 8197
rect 6010 8186 6016 8188
rect 6072 8186 6096 8188
rect 6152 8186 6176 8188
rect 6232 8186 6256 8188
rect 6312 8186 6318 8188
rect 6072 8134 6074 8186
rect 6254 8134 6256 8186
rect 6010 8132 6016 8134
rect 6072 8132 6096 8134
rect 6152 8132 6176 8134
rect 6232 8132 6256 8134
rect 6312 8132 6318 8134
rect 6010 8123 6318 8132
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5828 7546 5856 7822
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5816 7540 5868 7546
rect 5816 7482 5868 7488
rect 5920 7410 5948 7822
rect 6380 7410 6408 8434
rect 6670 7644 6978 7653
rect 6670 7642 6676 7644
rect 6732 7642 6756 7644
rect 6812 7642 6836 7644
rect 6892 7642 6916 7644
rect 6972 7642 6978 7644
rect 6732 7590 6734 7642
rect 6914 7590 6916 7642
rect 6670 7588 6676 7590
rect 6732 7588 6756 7590
rect 6812 7588 6836 7590
rect 6892 7588 6916 7590
rect 6972 7588 6978 7590
rect 6670 7579 6978 7588
rect 7760 7546 7788 8978
rect 8680 8945 8708 9046
rect 8666 8936 8722 8945
rect 8666 8871 8722 8880
rect 8694 8732 9002 8741
rect 8694 8730 8700 8732
rect 8756 8730 8780 8732
rect 8836 8730 8860 8732
rect 8916 8730 8940 8732
rect 8996 8730 9002 8732
rect 8756 8678 8758 8730
rect 8938 8678 8940 8730
rect 8694 8676 8700 8678
rect 8756 8676 8780 8678
rect 8836 8676 8860 8678
rect 8916 8676 8940 8678
rect 8996 8676 9002 8678
rect 8694 8667 9002 8676
rect 7932 8288 7984 8294
rect 7932 8230 7984 8236
rect 7944 7546 7972 8230
rect 8034 8188 8342 8197
rect 8034 8186 8040 8188
rect 8096 8186 8120 8188
rect 8176 8186 8200 8188
rect 8256 8186 8280 8188
rect 8336 8186 8342 8188
rect 8096 8134 8098 8186
rect 8278 8134 8280 8186
rect 8034 8132 8040 8134
rect 8096 8132 8120 8134
rect 8176 8132 8200 8134
rect 8256 8132 8280 8134
rect 8336 8132 8342 8134
rect 8034 8123 8342 8132
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 7748 7540 7800 7546
rect 7748 7482 7800 7488
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5632 7200 5684 7206
rect 5552 7148 5632 7154
rect 5552 7142 5684 7148
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 5460 7002 5488 7142
rect 5552 7126 5672 7142
rect 5448 6996 5500 7002
rect 5448 6938 5500 6944
rect 5356 6928 5408 6934
rect 5356 6870 5408 6876
rect 5172 6452 5224 6458
rect 5172 6394 5224 6400
rect 5080 5908 5132 5914
rect 5080 5850 5132 5856
rect 3884 5228 3936 5234
rect 3884 5170 3936 5176
rect 4356 5222 4476 5250
rect 4908 5222 5028 5250
rect 3986 4924 4294 4933
rect 3986 4922 3992 4924
rect 4048 4922 4072 4924
rect 4128 4922 4152 4924
rect 4208 4922 4232 4924
rect 4288 4922 4294 4924
rect 4048 4870 4050 4922
rect 4230 4870 4232 4922
rect 3986 4868 3992 4870
rect 4048 4868 4072 4870
rect 4128 4868 4152 4870
rect 4208 4868 4232 4870
rect 4288 4868 4294 4870
rect 3986 4859 4294 4868
rect 3608 4820 3660 4826
rect 3608 4762 3660 4768
rect 4356 4622 4384 5222
rect 4436 5160 4488 5166
rect 4436 5102 4488 5108
rect 3976 4616 4028 4622
rect 4344 4616 4396 4622
rect 3976 4558 4028 4564
rect 4264 4564 4344 4570
rect 4264 4558 4396 4564
rect 3988 4486 4016 4558
rect 4264 4542 4384 4558
rect 3148 4480 3200 4486
rect 3148 4422 3200 4428
rect 3516 4480 3568 4486
rect 3516 4422 3568 4428
rect 3976 4480 4028 4486
rect 3976 4422 4028 4428
rect 3056 4276 3108 4282
rect 3056 4218 3108 4224
rect 2964 3936 3016 3942
rect 2964 3878 3016 3884
rect 2622 3292 2930 3301
rect 2622 3290 2628 3292
rect 2684 3290 2708 3292
rect 2764 3290 2788 3292
rect 2844 3290 2868 3292
rect 2924 3290 2930 3292
rect 2684 3238 2686 3290
rect 2866 3238 2868 3290
rect 2622 3236 2628 3238
rect 2684 3236 2708 3238
rect 2764 3236 2788 3238
rect 2844 3236 2868 3238
rect 2924 3236 2930 3238
rect 2622 3227 2930 3236
rect 3160 3194 3188 4422
rect 4264 4282 4292 4542
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4252 4276 4304 4282
rect 4252 4218 4304 4224
rect 3986 3836 4294 3845
rect 3986 3834 3992 3836
rect 4048 3834 4072 3836
rect 4128 3834 4152 3836
rect 4208 3834 4232 3836
rect 4288 3834 4294 3836
rect 4048 3782 4050 3834
rect 4230 3782 4232 3834
rect 3986 3780 3992 3782
rect 4048 3780 4072 3782
rect 4128 3780 4152 3782
rect 4208 3780 4232 3782
rect 4288 3780 4294 3782
rect 3986 3771 4294 3780
rect 4252 3664 4304 3670
rect 4356 3618 4384 4422
rect 4304 3612 4384 3618
rect 4252 3606 4384 3612
rect 4264 3590 4384 3606
rect 3976 3460 4028 3466
rect 3976 3402 4028 3408
rect 3988 3346 4016 3402
rect 3896 3318 4016 3346
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 2596 3120 2648 3126
rect 2596 3062 2648 3068
rect 2608 2650 2636 3062
rect 3896 2666 3924 3318
rect 4264 2922 4292 3590
rect 4344 3392 4396 3398
rect 4344 3334 4396 3340
rect 4252 2916 4304 2922
rect 4252 2858 4304 2864
rect 3986 2748 4294 2757
rect 3986 2746 3992 2748
rect 4048 2746 4072 2748
rect 4128 2746 4152 2748
rect 4208 2746 4232 2748
rect 4288 2746 4294 2748
rect 4048 2694 4050 2746
rect 4230 2694 4232 2746
rect 3986 2692 3992 2694
rect 4048 2692 4072 2694
rect 4128 2692 4152 2694
rect 4208 2692 4232 2694
rect 4288 2692 4294 2694
rect 3986 2683 4294 2692
rect 3804 2650 3924 2666
rect 4356 2650 4384 3334
rect 4448 3058 4476 5102
rect 4712 5024 4764 5030
rect 4712 4966 4764 4972
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 4540 4162 4568 4762
rect 4724 4622 4752 4966
rect 4908 4622 4936 5222
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4896 4616 4948 4622
rect 4896 4558 4948 4564
rect 4988 4548 5040 4554
rect 4988 4490 5040 4496
rect 4646 4380 4954 4389
rect 4646 4378 4652 4380
rect 4708 4378 4732 4380
rect 4788 4378 4812 4380
rect 4868 4378 4892 4380
rect 4948 4378 4954 4380
rect 4708 4326 4710 4378
rect 4890 4326 4892 4378
rect 4646 4324 4652 4326
rect 4708 4324 4732 4326
rect 4788 4324 4812 4326
rect 4868 4324 4892 4326
rect 4948 4324 4954 4326
rect 4646 4315 4954 4324
rect 4712 4276 4764 4282
rect 4712 4218 4764 4224
rect 4540 4134 4660 4162
rect 4528 4072 4580 4078
rect 4528 4014 4580 4020
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 4436 2916 4488 2922
rect 4436 2858 4488 2864
rect 2596 2644 2648 2650
rect 2596 2586 2648 2592
rect 3792 2644 3924 2650
rect 3844 2638 3924 2644
rect 4344 2644 4396 2650
rect 3792 2586 3844 2592
rect 4344 2586 4396 2592
rect 2516 2502 2636 2530
rect 2608 2378 2636 2502
rect 4448 2446 4476 2858
rect 4540 2650 4568 4014
rect 4632 3738 4660 4134
rect 4620 3732 4672 3738
rect 4620 3674 4672 3680
rect 4724 3602 4752 4218
rect 5000 4026 5028 4490
rect 4908 3998 5028 4026
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4908 3398 4936 3998
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4896 3392 4948 3398
rect 4896 3334 4948 3340
rect 4646 3292 4954 3301
rect 4646 3290 4652 3292
rect 4708 3290 4732 3292
rect 4788 3290 4812 3292
rect 4868 3290 4892 3292
rect 4948 3290 4954 3292
rect 4708 3238 4710 3290
rect 4890 3238 4892 3290
rect 4646 3236 4652 3238
rect 4708 3236 4732 3238
rect 4788 3236 4812 3238
rect 4868 3236 4892 3238
rect 4948 3236 4954 3238
rect 4646 3227 4954 3236
rect 5000 3058 5028 3878
rect 5092 3126 5120 5850
rect 5184 5386 5212 6394
rect 5828 6322 5856 7142
rect 5920 6730 5948 7346
rect 6012 7206 6040 7346
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6010 7100 6318 7109
rect 6010 7098 6016 7100
rect 6072 7098 6096 7100
rect 6152 7098 6176 7100
rect 6232 7098 6256 7100
rect 6312 7098 6318 7100
rect 6072 7046 6074 7098
rect 6254 7046 6256 7098
rect 6010 7044 6016 7046
rect 6072 7044 6096 7046
rect 6152 7044 6176 7046
rect 6232 7044 6256 7046
rect 6312 7044 6318 7046
rect 6010 7035 6318 7044
rect 6380 6798 6408 7346
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 5908 6724 5960 6730
rect 5908 6666 5960 6672
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 6010 6012 6318 6021
rect 6010 6010 6016 6012
rect 6072 6010 6096 6012
rect 6152 6010 6176 6012
rect 6232 6010 6256 6012
rect 6312 6010 6318 6012
rect 6072 5958 6074 6010
rect 6254 5958 6256 6010
rect 6010 5956 6016 5958
rect 6072 5956 6096 5958
rect 6152 5956 6176 5958
rect 6232 5956 6256 5958
rect 6312 5956 6318 5958
rect 6010 5947 6318 5956
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 5632 5568 5684 5574
rect 5632 5510 5684 5516
rect 5184 5370 5304 5386
rect 5172 5364 5304 5370
rect 5224 5358 5304 5364
rect 5172 5306 5224 5312
rect 5172 5228 5224 5234
rect 5172 5170 5224 5176
rect 5184 4826 5212 5170
rect 5172 4820 5224 4826
rect 5172 4762 5224 4768
rect 5276 4706 5304 5358
rect 5184 4678 5396 4706
rect 5184 4282 5212 4678
rect 5172 4276 5224 4282
rect 5172 4218 5224 4224
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5184 3738 5212 3878
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5080 3120 5132 3126
rect 5080 3062 5132 3068
rect 4988 3052 5040 3058
rect 4988 2994 5040 3000
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 5184 2446 5212 3674
rect 5368 2446 5396 4678
rect 5644 4486 5672 5510
rect 6196 5234 6224 5646
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 6380 5166 6408 6734
rect 7392 6730 7420 7346
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7472 6928 7524 6934
rect 7472 6870 7524 6876
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 6670 6556 6978 6565
rect 6670 6554 6676 6556
rect 6732 6554 6756 6556
rect 6812 6554 6836 6556
rect 6892 6554 6916 6556
rect 6972 6554 6978 6556
rect 6732 6502 6734 6554
rect 6914 6502 6916 6554
rect 6670 6500 6676 6502
rect 6732 6500 6756 6502
rect 6812 6500 6836 6502
rect 6892 6500 6916 6502
rect 6972 6500 6978 6502
rect 6670 6491 6978 6500
rect 7392 6254 7420 6666
rect 7484 6458 7512 6870
rect 7656 6724 7708 6730
rect 7760 6712 7788 7142
rect 7944 6798 7972 7482
rect 8392 7268 8444 7274
rect 8392 7210 8444 7216
rect 8034 7100 8342 7109
rect 8034 7098 8040 7100
rect 8096 7098 8120 7100
rect 8176 7098 8200 7100
rect 8256 7098 8280 7100
rect 8336 7098 8342 7100
rect 8096 7046 8098 7098
rect 8278 7046 8280 7098
rect 8034 7044 8040 7046
rect 8096 7044 8120 7046
rect 8176 7044 8200 7046
rect 8256 7044 8280 7046
rect 8336 7044 8342 7046
rect 8034 7035 8342 7044
rect 7932 6792 7984 6798
rect 7932 6734 7984 6740
rect 7708 6684 7788 6712
rect 7656 6666 7708 6672
rect 7472 6452 7524 6458
rect 7472 6394 7524 6400
rect 7380 6248 7432 6254
rect 7380 6190 7432 6196
rect 7760 6202 7788 6684
rect 8404 6662 8432 7210
rect 8496 7002 8524 7822
rect 9128 7744 9180 7750
rect 9128 7686 9180 7692
rect 8694 7644 9002 7653
rect 8694 7642 8700 7644
rect 8756 7642 8780 7644
rect 8836 7642 8860 7644
rect 8916 7642 8940 7644
rect 8996 7642 9002 7644
rect 8756 7590 8758 7642
rect 8938 7590 8940 7642
rect 8694 7588 8700 7590
rect 8756 7588 8780 7590
rect 8836 7588 8860 7590
rect 8916 7588 8940 7590
rect 8996 7588 9002 7590
rect 8694 7579 9002 7588
rect 9140 7585 9168 7686
rect 9126 7576 9182 7585
rect 9126 7511 9182 7520
rect 8484 6996 8536 7002
rect 8484 6938 8536 6944
rect 8574 6896 8630 6905
rect 8574 6831 8576 6840
rect 8628 6831 8630 6840
rect 8576 6802 8628 6808
rect 8484 6792 8536 6798
rect 8484 6734 8536 6740
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 6474 8432 6598
rect 8312 6446 8432 6474
rect 8312 6390 8340 6446
rect 8300 6384 8352 6390
rect 8300 6326 8352 6332
rect 8496 6254 8524 6734
rect 8694 6556 9002 6565
rect 8694 6554 8700 6556
rect 8756 6554 8780 6556
rect 8836 6554 8860 6556
rect 8916 6554 8940 6556
rect 8996 6554 9002 6556
rect 8756 6502 8758 6554
rect 8938 6502 8940 6554
rect 8694 6500 8700 6502
rect 8756 6500 8780 6502
rect 8836 6500 8860 6502
rect 8916 6500 8940 6502
rect 8996 6500 9002 6502
rect 8694 6491 9002 6500
rect 8484 6248 8536 6254
rect 7760 6174 8064 6202
rect 8484 6190 8536 6196
rect 8666 6216 8722 6225
rect 8036 6118 8064 6174
rect 8666 6151 8722 6160
rect 7840 6112 7892 6118
rect 7840 6054 7892 6060
rect 7932 6112 7984 6118
rect 7932 6054 7984 6060
rect 8024 6112 8076 6118
rect 8024 6054 8076 6060
rect 7852 5794 7880 6054
rect 7944 5914 7972 6054
rect 8034 6012 8342 6021
rect 8034 6010 8040 6012
rect 8096 6010 8120 6012
rect 8176 6010 8200 6012
rect 8256 6010 8280 6012
rect 8336 6010 8342 6012
rect 8096 5958 8098 6010
rect 8278 5958 8280 6010
rect 8034 5956 8040 5958
rect 8096 5956 8120 5958
rect 8176 5956 8200 5958
rect 8256 5956 8280 5958
rect 8336 5956 8342 5958
rect 8034 5947 8342 5956
rect 8680 5914 8708 6151
rect 7932 5908 7984 5914
rect 7932 5850 7984 5856
rect 8668 5908 8720 5914
rect 8668 5850 8720 5856
rect 7852 5766 7972 5794
rect 7656 5704 7708 5710
rect 7656 5646 7708 5652
rect 6670 5468 6978 5477
rect 6670 5466 6676 5468
rect 6732 5466 6756 5468
rect 6812 5466 6836 5468
rect 6892 5466 6916 5468
rect 6972 5466 6978 5468
rect 6732 5414 6734 5466
rect 6914 5414 6916 5466
rect 6670 5412 6676 5414
rect 6732 5412 6756 5414
rect 6812 5412 6836 5414
rect 6892 5412 6916 5414
rect 6972 5412 6978 5414
rect 6670 5403 6978 5412
rect 7472 5228 7524 5234
rect 7472 5170 7524 5176
rect 6368 5160 6420 5166
rect 6368 5102 6420 5108
rect 6010 4924 6318 4933
rect 6010 4922 6016 4924
rect 6072 4922 6096 4924
rect 6152 4922 6176 4924
rect 6232 4922 6256 4924
rect 6312 4922 6318 4924
rect 6072 4870 6074 4922
rect 6254 4870 6256 4922
rect 6010 4868 6016 4870
rect 6072 4868 6096 4870
rect 6152 4868 6176 4870
rect 6232 4868 6256 4870
rect 6312 4868 6318 4870
rect 6010 4859 6318 4868
rect 6380 4622 6408 5102
rect 7484 4758 7512 5170
rect 7668 4826 7696 5646
rect 7944 5642 7972 5766
rect 7932 5636 7984 5642
rect 7932 5578 7984 5584
rect 7840 5160 7892 5166
rect 7840 5102 7892 5108
rect 7748 5024 7800 5030
rect 7748 4966 7800 4972
rect 7656 4820 7708 4826
rect 7656 4762 7708 4768
rect 7472 4752 7524 4758
rect 7472 4694 7524 4700
rect 6368 4616 6420 4622
rect 6368 4558 6420 4564
rect 5632 4480 5684 4486
rect 5632 4422 5684 4428
rect 6010 3836 6318 3845
rect 6010 3834 6016 3836
rect 6072 3834 6096 3836
rect 6152 3834 6176 3836
rect 6232 3834 6256 3836
rect 6312 3834 6318 3836
rect 6072 3782 6074 3834
rect 6254 3782 6256 3834
rect 6010 3780 6016 3782
rect 6072 3780 6096 3782
rect 6152 3780 6176 3782
rect 6232 3780 6256 3782
rect 6312 3780 6318 3782
rect 6010 3771 6318 3780
rect 5448 3596 5500 3602
rect 5448 3538 5500 3544
rect 5460 3194 5488 3538
rect 6380 3466 6408 4558
rect 6670 4380 6978 4389
rect 6670 4378 6676 4380
rect 6732 4378 6756 4380
rect 6812 4378 6836 4380
rect 6892 4378 6916 4380
rect 6972 4378 6978 4380
rect 6732 4326 6734 4378
rect 6914 4326 6916 4378
rect 6670 4324 6676 4326
rect 6732 4324 6756 4326
rect 6812 4324 6836 4326
rect 6892 4324 6916 4326
rect 6972 4324 6978 4326
rect 6670 4315 6978 4324
rect 7484 4162 7512 4694
rect 7760 4622 7788 4966
rect 7852 4622 7880 5102
rect 7748 4616 7800 4622
rect 7748 4558 7800 4564
rect 7840 4616 7892 4622
rect 7840 4558 7892 4564
rect 7760 4282 7788 4558
rect 7748 4276 7800 4282
rect 7748 4218 7800 4224
rect 7484 4146 7604 4162
rect 7484 4140 7616 4146
rect 7484 4134 7564 4140
rect 7564 4082 7616 4088
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7656 3936 7708 3942
rect 7656 3878 7708 3884
rect 7668 3534 7696 3878
rect 7760 3738 7788 4082
rect 7748 3732 7800 3738
rect 7748 3674 7800 3680
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 6368 3460 6420 3466
rect 6368 3402 6420 3408
rect 5448 3188 5500 3194
rect 5448 3130 5500 3136
rect 6380 3058 6408 3402
rect 6670 3292 6978 3301
rect 6670 3290 6676 3292
rect 6732 3290 6756 3292
rect 6812 3290 6836 3292
rect 6892 3290 6916 3292
rect 6972 3290 6978 3292
rect 6732 3238 6734 3290
rect 6914 3238 6916 3290
rect 6670 3236 6676 3238
rect 6732 3236 6756 3238
rect 6812 3236 6836 3238
rect 6892 3236 6916 3238
rect 6972 3236 6978 3238
rect 6670 3227 6978 3236
rect 7668 3074 7696 3470
rect 7760 3194 7788 3674
rect 7852 3398 7880 4558
rect 7944 4078 7972 5578
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8312 5234 8340 5510
rect 8694 5468 9002 5477
rect 8694 5466 8700 5468
rect 8756 5466 8780 5468
rect 8836 5466 8860 5468
rect 8916 5466 8940 5468
rect 8996 5466 9002 5468
rect 8756 5414 8758 5466
rect 8938 5414 8940 5466
rect 8694 5412 8700 5414
rect 8756 5412 8780 5414
rect 8836 5412 8860 5414
rect 8916 5412 8940 5414
rect 8996 5412 9002 5414
rect 8694 5403 9002 5412
rect 8300 5228 8352 5234
rect 8300 5170 8352 5176
rect 8392 5024 8444 5030
rect 8392 4966 8444 4972
rect 8760 5024 8812 5030
rect 8760 4966 8812 4972
rect 8034 4924 8342 4933
rect 8034 4922 8040 4924
rect 8096 4922 8120 4924
rect 8176 4922 8200 4924
rect 8256 4922 8280 4924
rect 8336 4922 8342 4924
rect 8096 4870 8098 4922
rect 8278 4870 8280 4922
rect 8034 4868 8040 4870
rect 8096 4868 8120 4870
rect 8176 4868 8200 4870
rect 8256 4868 8280 4870
rect 8336 4868 8342 4870
rect 8034 4859 8342 4868
rect 8404 4826 8432 4966
rect 8772 4865 8800 4966
rect 8758 4856 8814 4865
rect 8392 4820 8444 4826
rect 8758 4791 8814 4800
rect 8392 4762 8444 4768
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 8694 4380 9002 4389
rect 8694 4378 8700 4380
rect 8756 4378 8780 4380
rect 8836 4378 8860 4380
rect 8916 4378 8940 4380
rect 8996 4378 9002 4380
rect 8756 4326 8758 4378
rect 8938 4326 8940 4378
rect 8694 4324 8700 4326
rect 8756 4324 8780 4326
rect 8836 4324 8860 4326
rect 8916 4324 8940 4326
rect 8996 4324 9002 4326
rect 8694 4315 9002 4324
rect 9140 4185 9168 4422
rect 9126 4176 9182 4185
rect 9126 4111 9182 4120
rect 7932 4072 7984 4078
rect 7932 4014 7984 4020
rect 8034 3836 8342 3845
rect 8034 3834 8040 3836
rect 8096 3834 8120 3836
rect 8176 3834 8200 3836
rect 8256 3834 8280 3836
rect 8336 3834 8342 3836
rect 8096 3782 8098 3834
rect 8278 3782 8280 3834
rect 8034 3780 8040 3782
rect 8096 3780 8120 3782
rect 8176 3780 8200 3782
rect 8256 3780 8280 3782
rect 8336 3780 8342 3782
rect 8034 3771 8342 3780
rect 8668 3664 8720 3670
rect 8668 3606 8720 3612
rect 8208 3528 8260 3534
rect 8680 3505 8708 3606
rect 8208 3470 8260 3476
rect 8666 3496 8722 3505
rect 7840 3392 7892 3398
rect 7840 3334 7892 3340
rect 7748 3188 7800 3194
rect 7748 3130 7800 3136
rect 7852 3126 7880 3334
rect 7840 3120 7892 3126
rect 6368 3052 6420 3058
rect 7668 3046 7788 3074
rect 8220 3108 8248 3470
rect 8666 3431 8722 3440
rect 8694 3292 9002 3301
rect 8694 3290 8700 3292
rect 8756 3290 8780 3292
rect 8836 3290 8860 3292
rect 8916 3290 8940 3292
rect 8996 3290 9002 3292
rect 8756 3238 8758 3290
rect 8938 3238 8940 3290
rect 8694 3236 8700 3238
rect 8756 3236 8780 3238
rect 8836 3236 8860 3238
rect 8916 3236 8940 3238
rect 8996 3236 9002 3238
rect 8694 3227 9002 3236
rect 7840 3062 7892 3068
rect 7944 3080 8248 3108
rect 6368 2994 6420 3000
rect 7760 2990 7788 3046
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 6010 2748 6318 2757
rect 6010 2746 6016 2748
rect 6072 2746 6096 2748
rect 6152 2746 6176 2748
rect 6232 2746 6256 2748
rect 6312 2746 6318 2748
rect 6072 2694 6074 2746
rect 6254 2694 6256 2746
rect 6010 2692 6016 2694
rect 6072 2692 6096 2694
rect 6152 2692 6176 2694
rect 6232 2692 6256 2694
rect 6312 2692 6318 2694
rect 6010 2683 6318 2692
rect 7760 2514 7788 2926
rect 7840 2848 7892 2854
rect 7840 2790 7892 2796
rect 7748 2508 7800 2514
rect 7748 2450 7800 2456
rect 7852 2446 7880 2790
rect 7944 2650 7972 3080
rect 8758 2816 8814 2825
rect 8034 2748 8342 2757
rect 8758 2751 8814 2760
rect 8034 2746 8040 2748
rect 8096 2746 8120 2748
rect 8176 2746 8200 2748
rect 8256 2746 8280 2748
rect 8336 2746 8342 2748
rect 8096 2694 8098 2746
rect 8278 2694 8280 2746
rect 8034 2692 8040 2694
rect 8096 2692 8120 2694
rect 8176 2692 8200 2694
rect 8256 2692 8280 2694
rect 8336 2692 8342 2694
rect 8034 2683 8342 2692
rect 8772 2650 8800 2751
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 4436 2440 4488 2446
rect 4436 2382 4488 2388
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5356 2440 5408 2446
rect 5356 2382 5408 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 2596 2372 2648 2378
rect 2596 2314 2648 2320
rect 2622 2204 2930 2213
rect 2622 2202 2628 2204
rect 2684 2202 2708 2204
rect 2764 2202 2788 2204
rect 2844 2202 2868 2204
rect 2924 2202 2930 2204
rect 2684 2150 2686 2202
rect 2866 2150 2868 2202
rect 2622 2148 2628 2150
rect 2684 2148 2708 2150
rect 2764 2148 2788 2150
rect 2844 2148 2868 2150
rect 2924 2148 2930 2150
rect 2622 2139 2930 2148
rect 4646 2204 4954 2213
rect 4646 2202 4652 2204
rect 4708 2202 4732 2204
rect 4788 2202 4812 2204
rect 4868 2202 4892 2204
rect 4948 2202 4954 2204
rect 4708 2150 4710 2202
rect 4890 2150 4892 2202
rect 4646 2148 4652 2150
rect 4708 2148 4732 2150
rect 4788 2148 4812 2150
rect 4868 2148 4892 2150
rect 4948 2148 4954 2150
rect 4646 2139 4954 2148
rect 6670 2204 6978 2213
rect 6670 2202 6676 2204
rect 6732 2202 6756 2204
rect 6812 2202 6836 2204
rect 6892 2202 6916 2204
rect 6972 2202 6978 2204
rect 6732 2150 6734 2202
rect 6914 2150 6916 2202
rect 6670 2148 6676 2150
rect 6732 2148 6756 2150
rect 6812 2148 6836 2150
rect 6892 2148 6916 2150
rect 6972 2148 6978 2150
rect 6670 2139 6978 2148
rect 8694 2204 9002 2213
rect 8694 2202 8700 2204
rect 8756 2202 8780 2204
rect 8836 2202 8860 2204
rect 8916 2202 8940 2204
rect 8996 2202 9002 2204
rect 8756 2150 8758 2202
rect 8938 2150 8940 2202
rect 8694 2148 8700 2150
rect 8756 2148 8780 2150
rect 8836 2148 8860 2150
rect 8916 2148 8940 2150
rect 8996 2148 9002 2150
rect 8694 2139 9002 2148
<< via2 >>
rect 2628 9818 2684 9820
rect 2708 9818 2764 9820
rect 2788 9818 2844 9820
rect 2868 9818 2924 9820
rect 2628 9766 2674 9818
rect 2674 9766 2684 9818
rect 2708 9766 2738 9818
rect 2738 9766 2750 9818
rect 2750 9766 2764 9818
rect 2788 9766 2802 9818
rect 2802 9766 2814 9818
rect 2814 9766 2844 9818
rect 2868 9766 2878 9818
rect 2878 9766 2924 9818
rect 2628 9764 2684 9766
rect 2708 9764 2764 9766
rect 2788 9764 2844 9766
rect 2868 9764 2924 9766
rect 4652 9818 4708 9820
rect 4732 9818 4788 9820
rect 4812 9818 4868 9820
rect 4892 9818 4948 9820
rect 4652 9766 4698 9818
rect 4698 9766 4708 9818
rect 4732 9766 4762 9818
rect 4762 9766 4774 9818
rect 4774 9766 4788 9818
rect 4812 9766 4826 9818
rect 4826 9766 4838 9818
rect 4838 9766 4868 9818
rect 4892 9766 4902 9818
rect 4902 9766 4948 9818
rect 4652 9764 4708 9766
rect 4732 9764 4788 9766
rect 4812 9764 4868 9766
rect 4892 9764 4948 9766
rect 6676 9818 6732 9820
rect 6756 9818 6812 9820
rect 6836 9818 6892 9820
rect 6916 9818 6972 9820
rect 6676 9766 6722 9818
rect 6722 9766 6732 9818
rect 6756 9766 6786 9818
rect 6786 9766 6798 9818
rect 6798 9766 6812 9818
rect 6836 9766 6850 9818
rect 6850 9766 6862 9818
rect 6862 9766 6892 9818
rect 6916 9766 6926 9818
rect 6926 9766 6972 9818
rect 6676 9764 6732 9766
rect 6756 9764 6812 9766
rect 6836 9764 6892 9766
rect 6916 9764 6972 9766
rect 8700 9818 8756 9820
rect 8780 9818 8836 9820
rect 8860 9818 8916 9820
rect 8940 9818 8996 9820
rect 8700 9766 8746 9818
rect 8746 9766 8756 9818
rect 8780 9766 8810 9818
rect 8810 9766 8822 9818
rect 8822 9766 8836 9818
rect 8860 9766 8874 9818
rect 8874 9766 8886 9818
rect 8886 9766 8916 9818
rect 8940 9766 8950 9818
rect 8950 9766 8996 9818
rect 8700 9764 8756 9766
rect 8780 9764 8836 9766
rect 8860 9764 8916 9766
rect 8940 9764 8996 9766
rect 1968 9274 2024 9276
rect 2048 9274 2104 9276
rect 2128 9274 2184 9276
rect 2208 9274 2264 9276
rect 1968 9222 2014 9274
rect 2014 9222 2024 9274
rect 2048 9222 2078 9274
rect 2078 9222 2090 9274
rect 2090 9222 2104 9274
rect 2128 9222 2142 9274
rect 2142 9222 2154 9274
rect 2154 9222 2184 9274
rect 2208 9222 2218 9274
rect 2218 9222 2264 9274
rect 1968 9220 2024 9222
rect 2048 9220 2104 9222
rect 2128 9220 2184 9222
rect 2208 9220 2264 9222
rect 3992 9274 4048 9276
rect 4072 9274 4128 9276
rect 4152 9274 4208 9276
rect 4232 9274 4288 9276
rect 3992 9222 4038 9274
rect 4038 9222 4048 9274
rect 4072 9222 4102 9274
rect 4102 9222 4114 9274
rect 4114 9222 4128 9274
rect 4152 9222 4166 9274
rect 4166 9222 4178 9274
rect 4178 9222 4208 9274
rect 4232 9222 4242 9274
rect 4242 9222 4288 9274
rect 3992 9220 4048 9222
rect 4072 9220 4128 9222
rect 4152 9220 4208 9222
rect 4232 9220 4288 9222
rect 6016 9274 6072 9276
rect 6096 9274 6152 9276
rect 6176 9274 6232 9276
rect 6256 9274 6312 9276
rect 6016 9222 6062 9274
rect 6062 9222 6072 9274
rect 6096 9222 6126 9274
rect 6126 9222 6138 9274
rect 6138 9222 6152 9274
rect 6176 9222 6190 9274
rect 6190 9222 6202 9274
rect 6202 9222 6232 9274
rect 6256 9222 6266 9274
rect 6266 9222 6312 9274
rect 6016 9220 6072 9222
rect 6096 9220 6152 9222
rect 6176 9220 6232 9222
rect 6256 9220 6312 9222
rect 8040 9274 8096 9276
rect 8120 9274 8176 9276
rect 8200 9274 8256 9276
rect 8280 9274 8336 9276
rect 8040 9222 8086 9274
rect 8086 9222 8096 9274
rect 8120 9222 8150 9274
rect 8150 9222 8162 9274
rect 8162 9222 8176 9274
rect 8200 9222 8214 9274
rect 8214 9222 8226 9274
rect 8226 9222 8256 9274
rect 8280 9222 8290 9274
rect 8290 9222 8336 9274
rect 8040 9220 8096 9222
rect 8120 9220 8176 9222
rect 8200 9220 8256 9222
rect 8280 9220 8336 9222
rect 3790 8880 3846 8936
rect 2628 8730 2684 8732
rect 2708 8730 2764 8732
rect 2788 8730 2844 8732
rect 2868 8730 2924 8732
rect 2628 8678 2674 8730
rect 2674 8678 2684 8730
rect 2708 8678 2738 8730
rect 2738 8678 2750 8730
rect 2750 8678 2764 8730
rect 2788 8678 2802 8730
rect 2802 8678 2814 8730
rect 2814 8678 2844 8730
rect 2868 8678 2878 8730
rect 2878 8678 2924 8730
rect 2628 8676 2684 8678
rect 2708 8676 2764 8678
rect 2788 8676 2844 8678
rect 2868 8676 2924 8678
rect 1968 8186 2024 8188
rect 2048 8186 2104 8188
rect 2128 8186 2184 8188
rect 2208 8186 2264 8188
rect 1968 8134 2014 8186
rect 2014 8134 2024 8186
rect 2048 8134 2078 8186
rect 2078 8134 2090 8186
rect 2090 8134 2104 8186
rect 2128 8134 2142 8186
rect 2142 8134 2154 8186
rect 2154 8134 2184 8186
rect 2208 8134 2218 8186
rect 2218 8134 2264 8186
rect 1968 8132 2024 8134
rect 2048 8132 2104 8134
rect 2128 8132 2184 8134
rect 2208 8132 2264 8134
rect 1398 7520 1454 7576
rect 2628 7642 2684 7644
rect 2708 7642 2764 7644
rect 2788 7642 2844 7644
rect 2868 7642 2924 7644
rect 2628 7590 2674 7642
rect 2674 7590 2684 7642
rect 2708 7590 2738 7642
rect 2738 7590 2750 7642
rect 2750 7590 2764 7642
rect 2788 7590 2802 7642
rect 2802 7590 2814 7642
rect 2814 7590 2844 7642
rect 2868 7590 2878 7642
rect 2878 7590 2924 7642
rect 2628 7588 2684 7590
rect 2708 7588 2764 7590
rect 2788 7588 2844 7590
rect 2868 7588 2924 7590
rect 3514 7828 3516 7848
rect 3516 7828 3568 7848
rect 3568 7828 3570 7848
rect 3514 7792 3570 7828
rect 1968 7098 2024 7100
rect 2048 7098 2104 7100
rect 2128 7098 2184 7100
rect 2208 7098 2264 7100
rect 1968 7046 2014 7098
rect 2014 7046 2024 7098
rect 2048 7046 2078 7098
rect 2078 7046 2090 7098
rect 2090 7046 2104 7098
rect 2128 7046 2142 7098
rect 2142 7046 2154 7098
rect 2154 7046 2184 7098
rect 2208 7046 2218 7098
rect 2218 7046 2264 7098
rect 1968 7044 2024 7046
rect 2048 7044 2104 7046
rect 2128 7044 2184 7046
rect 2208 7044 2264 7046
rect 754 5908 810 5944
rect 754 5888 756 5908
rect 756 5888 808 5908
rect 808 5888 810 5908
rect 1968 6010 2024 6012
rect 2048 6010 2104 6012
rect 2128 6010 2184 6012
rect 2208 6010 2264 6012
rect 1968 5958 2014 6010
rect 2014 5958 2024 6010
rect 2048 5958 2078 6010
rect 2078 5958 2090 6010
rect 2090 5958 2104 6010
rect 2128 5958 2142 6010
rect 2142 5958 2154 6010
rect 2154 5958 2184 6010
rect 2208 5958 2218 6010
rect 2218 5958 2264 6010
rect 1968 5956 2024 5958
rect 2048 5956 2104 5958
rect 2128 5956 2184 5958
rect 2208 5956 2264 5958
rect 2628 6554 2684 6556
rect 2708 6554 2764 6556
rect 2788 6554 2844 6556
rect 2868 6554 2924 6556
rect 2628 6502 2674 6554
rect 2674 6502 2684 6554
rect 2708 6502 2738 6554
rect 2738 6502 2750 6554
rect 2750 6502 2764 6554
rect 2788 6502 2802 6554
rect 2802 6502 2814 6554
rect 2814 6502 2844 6554
rect 2868 6502 2878 6554
rect 2878 6502 2924 6554
rect 2628 6500 2684 6502
rect 2708 6500 2764 6502
rect 2788 6500 2844 6502
rect 2868 6500 2924 6502
rect 2628 5466 2684 5468
rect 2708 5466 2764 5468
rect 2788 5466 2844 5468
rect 2868 5466 2924 5468
rect 2628 5414 2674 5466
rect 2674 5414 2684 5466
rect 2708 5414 2738 5466
rect 2738 5414 2750 5466
rect 2750 5414 2764 5466
rect 2788 5414 2802 5466
rect 2802 5414 2814 5466
rect 2814 5414 2844 5466
rect 2868 5414 2878 5466
rect 2878 5414 2924 5466
rect 2628 5412 2684 5414
rect 2708 5412 2764 5414
rect 2788 5412 2844 5414
rect 2868 5412 2924 5414
rect 1968 4922 2024 4924
rect 2048 4922 2104 4924
rect 2128 4922 2184 4924
rect 2208 4922 2264 4924
rect 1968 4870 2014 4922
rect 2014 4870 2024 4922
rect 2048 4870 2078 4922
rect 2078 4870 2090 4922
rect 2090 4870 2104 4922
rect 2128 4870 2142 4922
rect 2142 4870 2154 4922
rect 2154 4870 2184 4922
rect 2208 4870 2218 4922
rect 2218 4870 2264 4922
rect 1968 4868 2024 4870
rect 2048 4868 2104 4870
rect 2128 4868 2184 4870
rect 2208 4868 2264 4870
rect 2628 4378 2684 4380
rect 2708 4378 2764 4380
rect 2788 4378 2844 4380
rect 2868 4378 2924 4380
rect 2628 4326 2674 4378
rect 2674 4326 2684 4378
rect 2708 4326 2738 4378
rect 2738 4326 2750 4378
rect 2750 4326 2764 4378
rect 2788 4326 2802 4378
rect 2802 4326 2814 4378
rect 2814 4326 2844 4378
rect 2868 4326 2878 4378
rect 2878 4326 2924 4378
rect 2628 4324 2684 4326
rect 2708 4324 2764 4326
rect 2788 4324 2844 4326
rect 2868 4324 2924 4326
rect 1968 3834 2024 3836
rect 2048 3834 2104 3836
rect 2128 3834 2184 3836
rect 2208 3834 2264 3836
rect 1968 3782 2014 3834
rect 2014 3782 2024 3834
rect 2048 3782 2078 3834
rect 2078 3782 2090 3834
rect 2090 3782 2104 3834
rect 2128 3782 2142 3834
rect 2142 3782 2154 3834
rect 2154 3782 2184 3834
rect 2208 3782 2218 3834
rect 2218 3782 2264 3834
rect 1968 3780 2024 3782
rect 2048 3780 2104 3782
rect 2128 3780 2184 3782
rect 2208 3780 2264 3782
rect 1968 2746 2024 2748
rect 2048 2746 2104 2748
rect 2128 2746 2184 2748
rect 2208 2746 2264 2748
rect 1968 2694 2014 2746
rect 2014 2694 2024 2746
rect 2048 2694 2078 2746
rect 2078 2694 2090 2746
rect 2090 2694 2104 2746
rect 2128 2694 2142 2746
rect 2142 2694 2154 2746
rect 2154 2694 2184 2746
rect 2208 2694 2218 2746
rect 2218 2694 2264 2746
rect 1968 2692 2024 2694
rect 2048 2692 2104 2694
rect 2128 2692 2184 2694
rect 2208 2692 2264 2694
rect 3992 8186 4048 8188
rect 4072 8186 4128 8188
rect 4152 8186 4208 8188
rect 4232 8186 4288 8188
rect 3992 8134 4038 8186
rect 4038 8134 4048 8186
rect 4072 8134 4102 8186
rect 4102 8134 4114 8186
rect 4114 8134 4128 8186
rect 4152 8134 4166 8186
rect 4166 8134 4178 8186
rect 4178 8134 4208 8186
rect 4232 8134 4242 8186
rect 4242 8134 4288 8186
rect 3992 8132 4048 8134
rect 4072 8132 4128 8134
rect 4152 8132 4208 8134
rect 4232 8132 4288 8134
rect 4652 8730 4708 8732
rect 4732 8730 4788 8732
rect 4812 8730 4868 8732
rect 4892 8730 4948 8732
rect 4652 8678 4698 8730
rect 4698 8678 4708 8730
rect 4732 8678 4762 8730
rect 4762 8678 4774 8730
rect 4774 8678 4788 8730
rect 4812 8678 4826 8730
rect 4826 8678 4838 8730
rect 4838 8678 4868 8730
rect 4892 8678 4902 8730
rect 4902 8678 4948 8730
rect 4652 8676 4708 8678
rect 4732 8676 4788 8678
rect 4812 8676 4868 8678
rect 4892 8676 4948 8678
rect 4434 7812 4490 7848
rect 4434 7792 4436 7812
rect 4436 7792 4488 7812
rect 4488 7792 4490 7812
rect 4652 7642 4708 7644
rect 4732 7642 4788 7644
rect 4812 7642 4868 7644
rect 4892 7642 4948 7644
rect 4652 7590 4698 7642
rect 4698 7590 4708 7642
rect 4732 7590 4762 7642
rect 4762 7590 4774 7642
rect 4774 7590 4788 7642
rect 4812 7590 4826 7642
rect 4826 7590 4838 7642
rect 4838 7590 4868 7642
rect 4892 7590 4902 7642
rect 4902 7590 4948 7642
rect 4652 7588 4708 7590
rect 4732 7588 4788 7590
rect 4812 7588 4868 7590
rect 4892 7588 4948 7590
rect 3992 7098 4048 7100
rect 4072 7098 4128 7100
rect 4152 7098 4208 7100
rect 4232 7098 4288 7100
rect 3992 7046 4038 7098
rect 4038 7046 4048 7098
rect 4072 7046 4102 7098
rect 4102 7046 4114 7098
rect 4114 7046 4128 7098
rect 4152 7046 4166 7098
rect 4166 7046 4178 7098
rect 4178 7046 4208 7098
rect 4232 7046 4242 7098
rect 4242 7046 4288 7098
rect 3992 7044 4048 7046
rect 4072 7044 4128 7046
rect 4152 7044 4208 7046
rect 4232 7044 4288 7046
rect 4652 6554 4708 6556
rect 4732 6554 4788 6556
rect 4812 6554 4868 6556
rect 4892 6554 4948 6556
rect 4652 6502 4698 6554
rect 4698 6502 4708 6554
rect 4732 6502 4762 6554
rect 4762 6502 4774 6554
rect 4774 6502 4788 6554
rect 4812 6502 4826 6554
rect 4826 6502 4838 6554
rect 4838 6502 4868 6554
rect 4892 6502 4902 6554
rect 4902 6502 4948 6554
rect 4652 6500 4708 6502
rect 4732 6500 4788 6502
rect 4812 6500 4868 6502
rect 4892 6500 4948 6502
rect 3992 6010 4048 6012
rect 4072 6010 4128 6012
rect 4152 6010 4208 6012
rect 4232 6010 4288 6012
rect 3992 5958 4038 6010
rect 4038 5958 4048 6010
rect 4072 5958 4102 6010
rect 4102 5958 4114 6010
rect 4114 5958 4128 6010
rect 4152 5958 4166 6010
rect 4166 5958 4178 6010
rect 4178 5958 4208 6010
rect 4232 5958 4242 6010
rect 4242 5958 4288 6010
rect 3992 5956 4048 5958
rect 4072 5956 4128 5958
rect 4152 5956 4208 5958
rect 4232 5956 4288 5958
rect 4652 5466 4708 5468
rect 4732 5466 4788 5468
rect 4812 5466 4868 5468
rect 4892 5466 4948 5468
rect 4652 5414 4698 5466
rect 4698 5414 4708 5466
rect 4732 5414 4762 5466
rect 4762 5414 4774 5466
rect 4774 5414 4788 5466
rect 4812 5414 4826 5466
rect 4826 5414 4838 5466
rect 4838 5414 4868 5466
rect 4892 5414 4902 5466
rect 4902 5414 4948 5466
rect 4652 5412 4708 5414
rect 4732 5412 4788 5414
rect 4812 5412 4868 5414
rect 4892 5412 4948 5414
rect 6676 8730 6732 8732
rect 6756 8730 6812 8732
rect 6836 8730 6892 8732
rect 6916 8730 6972 8732
rect 6676 8678 6722 8730
rect 6722 8678 6732 8730
rect 6756 8678 6786 8730
rect 6786 8678 6798 8730
rect 6798 8678 6812 8730
rect 6836 8678 6850 8730
rect 6850 8678 6862 8730
rect 6862 8678 6892 8730
rect 6916 8678 6926 8730
rect 6926 8678 6972 8730
rect 6676 8676 6732 8678
rect 6756 8676 6812 8678
rect 6836 8676 6892 8678
rect 6916 8676 6972 8678
rect 6016 8186 6072 8188
rect 6096 8186 6152 8188
rect 6176 8186 6232 8188
rect 6256 8186 6312 8188
rect 6016 8134 6062 8186
rect 6062 8134 6072 8186
rect 6096 8134 6126 8186
rect 6126 8134 6138 8186
rect 6138 8134 6152 8186
rect 6176 8134 6190 8186
rect 6190 8134 6202 8186
rect 6202 8134 6232 8186
rect 6256 8134 6266 8186
rect 6266 8134 6312 8186
rect 6016 8132 6072 8134
rect 6096 8132 6152 8134
rect 6176 8132 6232 8134
rect 6256 8132 6312 8134
rect 6676 7642 6732 7644
rect 6756 7642 6812 7644
rect 6836 7642 6892 7644
rect 6916 7642 6972 7644
rect 6676 7590 6722 7642
rect 6722 7590 6732 7642
rect 6756 7590 6786 7642
rect 6786 7590 6798 7642
rect 6798 7590 6812 7642
rect 6836 7590 6850 7642
rect 6850 7590 6862 7642
rect 6862 7590 6892 7642
rect 6916 7590 6926 7642
rect 6926 7590 6972 7642
rect 6676 7588 6732 7590
rect 6756 7588 6812 7590
rect 6836 7588 6892 7590
rect 6916 7588 6972 7590
rect 8666 8880 8722 8936
rect 8700 8730 8756 8732
rect 8780 8730 8836 8732
rect 8860 8730 8916 8732
rect 8940 8730 8996 8732
rect 8700 8678 8746 8730
rect 8746 8678 8756 8730
rect 8780 8678 8810 8730
rect 8810 8678 8822 8730
rect 8822 8678 8836 8730
rect 8860 8678 8874 8730
rect 8874 8678 8886 8730
rect 8886 8678 8916 8730
rect 8940 8678 8950 8730
rect 8950 8678 8996 8730
rect 8700 8676 8756 8678
rect 8780 8676 8836 8678
rect 8860 8676 8916 8678
rect 8940 8676 8996 8678
rect 8040 8186 8096 8188
rect 8120 8186 8176 8188
rect 8200 8186 8256 8188
rect 8280 8186 8336 8188
rect 8040 8134 8086 8186
rect 8086 8134 8096 8186
rect 8120 8134 8150 8186
rect 8150 8134 8162 8186
rect 8162 8134 8176 8186
rect 8200 8134 8214 8186
rect 8214 8134 8226 8186
rect 8226 8134 8256 8186
rect 8280 8134 8290 8186
rect 8290 8134 8336 8186
rect 8040 8132 8096 8134
rect 8120 8132 8176 8134
rect 8200 8132 8256 8134
rect 8280 8132 8336 8134
rect 3992 4922 4048 4924
rect 4072 4922 4128 4924
rect 4152 4922 4208 4924
rect 4232 4922 4288 4924
rect 3992 4870 4038 4922
rect 4038 4870 4048 4922
rect 4072 4870 4102 4922
rect 4102 4870 4114 4922
rect 4114 4870 4128 4922
rect 4152 4870 4166 4922
rect 4166 4870 4178 4922
rect 4178 4870 4208 4922
rect 4232 4870 4242 4922
rect 4242 4870 4288 4922
rect 3992 4868 4048 4870
rect 4072 4868 4128 4870
rect 4152 4868 4208 4870
rect 4232 4868 4288 4870
rect 2628 3290 2684 3292
rect 2708 3290 2764 3292
rect 2788 3290 2844 3292
rect 2868 3290 2924 3292
rect 2628 3238 2674 3290
rect 2674 3238 2684 3290
rect 2708 3238 2738 3290
rect 2738 3238 2750 3290
rect 2750 3238 2764 3290
rect 2788 3238 2802 3290
rect 2802 3238 2814 3290
rect 2814 3238 2844 3290
rect 2868 3238 2878 3290
rect 2878 3238 2924 3290
rect 2628 3236 2684 3238
rect 2708 3236 2764 3238
rect 2788 3236 2844 3238
rect 2868 3236 2924 3238
rect 3992 3834 4048 3836
rect 4072 3834 4128 3836
rect 4152 3834 4208 3836
rect 4232 3834 4288 3836
rect 3992 3782 4038 3834
rect 4038 3782 4048 3834
rect 4072 3782 4102 3834
rect 4102 3782 4114 3834
rect 4114 3782 4128 3834
rect 4152 3782 4166 3834
rect 4166 3782 4178 3834
rect 4178 3782 4208 3834
rect 4232 3782 4242 3834
rect 4242 3782 4288 3834
rect 3992 3780 4048 3782
rect 4072 3780 4128 3782
rect 4152 3780 4208 3782
rect 4232 3780 4288 3782
rect 3992 2746 4048 2748
rect 4072 2746 4128 2748
rect 4152 2746 4208 2748
rect 4232 2746 4288 2748
rect 3992 2694 4038 2746
rect 4038 2694 4048 2746
rect 4072 2694 4102 2746
rect 4102 2694 4114 2746
rect 4114 2694 4128 2746
rect 4152 2694 4166 2746
rect 4166 2694 4178 2746
rect 4178 2694 4208 2746
rect 4232 2694 4242 2746
rect 4242 2694 4288 2746
rect 3992 2692 4048 2694
rect 4072 2692 4128 2694
rect 4152 2692 4208 2694
rect 4232 2692 4288 2694
rect 4652 4378 4708 4380
rect 4732 4378 4788 4380
rect 4812 4378 4868 4380
rect 4892 4378 4948 4380
rect 4652 4326 4698 4378
rect 4698 4326 4708 4378
rect 4732 4326 4762 4378
rect 4762 4326 4774 4378
rect 4774 4326 4788 4378
rect 4812 4326 4826 4378
rect 4826 4326 4838 4378
rect 4838 4326 4868 4378
rect 4892 4326 4902 4378
rect 4902 4326 4948 4378
rect 4652 4324 4708 4326
rect 4732 4324 4788 4326
rect 4812 4324 4868 4326
rect 4892 4324 4948 4326
rect 4652 3290 4708 3292
rect 4732 3290 4788 3292
rect 4812 3290 4868 3292
rect 4892 3290 4948 3292
rect 4652 3238 4698 3290
rect 4698 3238 4708 3290
rect 4732 3238 4762 3290
rect 4762 3238 4774 3290
rect 4774 3238 4788 3290
rect 4812 3238 4826 3290
rect 4826 3238 4838 3290
rect 4838 3238 4868 3290
rect 4892 3238 4902 3290
rect 4902 3238 4948 3290
rect 4652 3236 4708 3238
rect 4732 3236 4788 3238
rect 4812 3236 4868 3238
rect 4892 3236 4948 3238
rect 6016 7098 6072 7100
rect 6096 7098 6152 7100
rect 6176 7098 6232 7100
rect 6256 7098 6312 7100
rect 6016 7046 6062 7098
rect 6062 7046 6072 7098
rect 6096 7046 6126 7098
rect 6126 7046 6138 7098
rect 6138 7046 6152 7098
rect 6176 7046 6190 7098
rect 6190 7046 6202 7098
rect 6202 7046 6232 7098
rect 6256 7046 6266 7098
rect 6266 7046 6312 7098
rect 6016 7044 6072 7046
rect 6096 7044 6152 7046
rect 6176 7044 6232 7046
rect 6256 7044 6312 7046
rect 6016 6010 6072 6012
rect 6096 6010 6152 6012
rect 6176 6010 6232 6012
rect 6256 6010 6312 6012
rect 6016 5958 6062 6010
rect 6062 5958 6072 6010
rect 6096 5958 6126 6010
rect 6126 5958 6138 6010
rect 6138 5958 6152 6010
rect 6176 5958 6190 6010
rect 6190 5958 6202 6010
rect 6202 5958 6232 6010
rect 6256 5958 6266 6010
rect 6266 5958 6312 6010
rect 6016 5956 6072 5958
rect 6096 5956 6152 5958
rect 6176 5956 6232 5958
rect 6256 5956 6312 5958
rect 6676 6554 6732 6556
rect 6756 6554 6812 6556
rect 6836 6554 6892 6556
rect 6916 6554 6972 6556
rect 6676 6502 6722 6554
rect 6722 6502 6732 6554
rect 6756 6502 6786 6554
rect 6786 6502 6798 6554
rect 6798 6502 6812 6554
rect 6836 6502 6850 6554
rect 6850 6502 6862 6554
rect 6862 6502 6892 6554
rect 6916 6502 6926 6554
rect 6926 6502 6972 6554
rect 6676 6500 6732 6502
rect 6756 6500 6812 6502
rect 6836 6500 6892 6502
rect 6916 6500 6972 6502
rect 8040 7098 8096 7100
rect 8120 7098 8176 7100
rect 8200 7098 8256 7100
rect 8280 7098 8336 7100
rect 8040 7046 8086 7098
rect 8086 7046 8096 7098
rect 8120 7046 8150 7098
rect 8150 7046 8162 7098
rect 8162 7046 8176 7098
rect 8200 7046 8214 7098
rect 8214 7046 8226 7098
rect 8226 7046 8256 7098
rect 8280 7046 8290 7098
rect 8290 7046 8336 7098
rect 8040 7044 8096 7046
rect 8120 7044 8176 7046
rect 8200 7044 8256 7046
rect 8280 7044 8336 7046
rect 8700 7642 8756 7644
rect 8780 7642 8836 7644
rect 8860 7642 8916 7644
rect 8940 7642 8996 7644
rect 8700 7590 8746 7642
rect 8746 7590 8756 7642
rect 8780 7590 8810 7642
rect 8810 7590 8822 7642
rect 8822 7590 8836 7642
rect 8860 7590 8874 7642
rect 8874 7590 8886 7642
rect 8886 7590 8916 7642
rect 8940 7590 8950 7642
rect 8950 7590 8996 7642
rect 8700 7588 8756 7590
rect 8780 7588 8836 7590
rect 8860 7588 8916 7590
rect 8940 7588 8996 7590
rect 9126 7520 9182 7576
rect 8574 6860 8630 6896
rect 8574 6840 8576 6860
rect 8576 6840 8628 6860
rect 8628 6840 8630 6860
rect 8700 6554 8756 6556
rect 8780 6554 8836 6556
rect 8860 6554 8916 6556
rect 8940 6554 8996 6556
rect 8700 6502 8746 6554
rect 8746 6502 8756 6554
rect 8780 6502 8810 6554
rect 8810 6502 8822 6554
rect 8822 6502 8836 6554
rect 8860 6502 8874 6554
rect 8874 6502 8886 6554
rect 8886 6502 8916 6554
rect 8940 6502 8950 6554
rect 8950 6502 8996 6554
rect 8700 6500 8756 6502
rect 8780 6500 8836 6502
rect 8860 6500 8916 6502
rect 8940 6500 8996 6502
rect 8666 6160 8722 6216
rect 8040 6010 8096 6012
rect 8120 6010 8176 6012
rect 8200 6010 8256 6012
rect 8280 6010 8336 6012
rect 8040 5958 8086 6010
rect 8086 5958 8096 6010
rect 8120 5958 8150 6010
rect 8150 5958 8162 6010
rect 8162 5958 8176 6010
rect 8200 5958 8214 6010
rect 8214 5958 8226 6010
rect 8226 5958 8256 6010
rect 8280 5958 8290 6010
rect 8290 5958 8336 6010
rect 8040 5956 8096 5958
rect 8120 5956 8176 5958
rect 8200 5956 8256 5958
rect 8280 5956 8336 5958
rect 6676 5466 6732 5468
rect 6756 5466 6812 5468
rect 6836 5466 6892 5468
rect 6916 5466 6972 5468
rect 6676 5414 6722 5466
rect 6722 5414 6732 5466
rect 6756 5414 6786 5466
rect 6786 5414 6798 5466
rect 6798 5414 6812 5466
rect 6836 5414 6850 5466
rect 6850 5414 6862 5466
rect 6862 5414 6892 5466
rect 6916 5414 6926 5466
rect 6926 5414 6972 5466
rect 6676 5412 6732 5414
rect 6756 5412 6812 5414
rect 6836 5412 6892 5414
rect 6916 5412 6972 5414
rect 6016 4922 6072 4924
rect 6096 4922 6152 4924
rect 6176 4922 6232 4924
rect 6256 4922 6312 4924
rect 6016 4870 6062 4922
rect 6062 4870 6072 4922
rect 6096 4870 6126 4922
rect 6126 4870 6138 4922
rect 6138 4870 6152 4922
rect 6176 4870 6190 4922
rect 6190 4870 6202 4922
rect 6202 4870 6232 4922
rect 6256 4870 6266 4922
rect 6266 4870 6312 4922
rect 6016 4868 6072 4870
rect 6096 4868 6152 4870
rect 6176 4868 6232 4870
rect 6256 4868 6312 4870
rect 6016 3834 6072 3836
rect 6096 3834 6152 3836
rect 6176 3834 6232 3836
rect 6256 3834 6312 3836
rect 6016 3782 6062 3834
rect 6062 3782 6072 3834
rect 6096 3782 6126 3834
rect 6126 3782 6138 3834
rect 6138 3782 6152 3834
rect 6176 3782 6190 3834
rect 6190 3782 6202 3834
rect 6202 3782 6232 3834
rect 6256 3782 6266 3834
rect 6266 3782 6312 3834
rect 6016 3780 6072 3782
rect 6096 3780 6152 3782
rect 6176 3780 6232 3782
rect 6256 3780 6312 3782
rect 6676 4378 6732 4380
rect 6756 4378 6812 4380
rect 6836 4378 6892 4380
rect 6916 4378 6972 4380
rect 6676 4326 6722 4378
rect 6722 4326 6732 4378
rect 6756 4326 6786 4378
rect 6786 4326 6798 4378
rect 6798 4326 6812 4378
rect 6836 4326 6850 4378
rect 6850 4326 6862 4378
rect 6862 4326 6892 4378
rect 6916 4326 6926 4378
rect 6926 4326 6972 4378
rect 6676 4324 6732 4326
rect 6756 4324 6812 4326
rect 6836 4324 6892 4326
rect 6916 4324 6972 4326
rect 6676 3290 6732 3292
rect 6756 3290 6812 3292
rect 6836 3290 6892 3292
rect 6916 3290 6972 3292
rect 6676 3238 6722 3290
rect 6722 3238 6732 3290
rect 6756 3238 6786 3290
rect 6786 3238 6798 3290
rect 6798 3238 6812 3290
rect 6836 3238 6850 3290
rect 6850 3238 6862 3290
rect 6862 3238 6892 3290
rect 6916 3238 6926 3290
rect 6926 3238 6972 3290
rect 6676 3236 6732 3238
rect 6756 3236 6812 3238
rect 6836 3236 6892 3238
rect 6916 3236 6972 3238
rect 8700 5466 8756 5468
rect 8780 5466 8836 5468
rect 8860 5466 8916 5468
rect 8940 5466 8996 5468
rect 8700 5414 8746 5466
rect 8746 5414 8756 5466
rect 8780 5414 8810 5466
rect 8810 5414 8822 5466
rect 8822 5414 8836 5466
rect 8860 5414 8874 5466
rect 8874 5414 8886 5466
rect 8886 5414 8916 5466
rect 8940 5414 8950 5466
rect 8950 5414 8996 5466
rect 8700 5412 8756 5414
rect 8780 5412 8836 5414
rect 8860 5412 8916 5414
rect 8940 5412 8996 5414
rect 8040 4922 8096 4924
rect 8120 4922 8176 4924
rect 8200 4922 8256 4924
rect 8280 4922 8336 4924
rect 8040 4870 8086 4922
rect 8086 4870 8096 4922
rect 8120 4870 8150 4922
rect 8150 4870 8162 4922
rect 8162 4870 8176 4922
rect 8200 4870 8214 4922
rect 8214 4870 8226 4922
rect 8226 4870 8256 4922
rect 8280 4870 8290 4922
rect 8290 4870 8336 4922
rect 8040 4868 8096 4870
rect 8120 4868 8176 4870
rect 8200 4868 8256 4870
rect 8280 4868 8336 4870
rect 8758 4800 8814 4856
rect 8700 4378 8756 4380
rect 8780 4378 8836 4380
rect 8860 4378 8916 4380
rect 8940 4378 8996 4380
rect 8700 4326 8746 4378
rect 8746 4326 8756 4378
rect 8780 4326 8810 4378
rect 8810 4326 8822 4378
rect 8822 4326 8836 4378
rect 8860 4326 8874 4378
rect 8874 4326 8886 4378
rect 8886 4326 8916 4378
rect 8940 4326 8950 4378
rect 8950 4326 8996 4378
rect 8700 4324 8756 4326
rect 8780 4324 8836 4326
rect 8860 4324 8916 4326
rect 8940 4324 8996 4326
rect 9126 4120 9182 4176
rect 8040 3834 8096 3836
rect 8120 3834 8176 3836
rect 8200 3834 8256 3836
rect 8280 3834 8336 3836
rect 8040 3782 8086 3834
rect 8086 3782 8096 3834
rect 8120 3782 8150 3834
rect 8150 3782 8162 3834
rect 8162 3782 8176 3834
rect 8200 3782 8214 3834
rect 8214 3782 8226 3834
rect 8226 3782 8256 3834
rect 8280 3782 8290 3834
rect 8290 3782 8336 3834
rect 8040 3780 8096 3782
rect 8120 3780 8176 3782
rect 8200 3780 8256 3782
rect 8280 3780 8336 3782
rect 8666 3440 8722 3496
rect 8700 3290 8756 3292
rect 8780 3290 8836 3292
rect 8860 3290 8916 3292
rect 8940 3290 8996 3292
rect 8700 3238 8746 3290
rect 8746 3238 8756 3290
rect 8780 3238 8810 3290
rect 8810 3238 8822 3290
rect 8822 3238 8836 3290
rect 8860 3238 8874 3290
rect 8874 3238 8886 3290
rect 8886 3238 8916 3290
rect 8940 3238 8950 3290
rect 8950 3238 8996 3290
rect 8700 3236 8756 3238
rect 8780 3236 8836 3238
rect 8860 3236 8916 3238
rect 8940 3236 8996 3238
rect 6016 2746 6072 2748
rect 6096 2746 6152 2748
rect 6176 2746 6232 2748
rect 6256 2746 6312 2748
rect 6016 2694 6062 2746
rect 6062 2694 6072 2746
rect 6096 2694 6126 2746
rect 6126 2694 6138 2746
rect 6138 2694 6152 2746
rect 6176 2694 6190 2746
rect 6190 2694 6202 2746
rect 6202 2694 6232 2746
rect 6256 2694 6266 2746
rect 6266 2694 6312 2746
rect 6016 2692 6072 2694
rect 6096 2692 6152 2694
rect 6176 2692 6232 2694
rect 6256 2692 6312 2694
rect 8758 2760 8814 2816
rect 8040 2746 8096 2748
rect 8120 2746 8176 2748
rect 8200 2746 8256 2748
rect 8280 2746 8336 2748
rect 8040 2694 8086 2746
rect 8086 2694 8096 2746
rect 8120 2694 8150 2746
rect 8150 2694 8162 2746
rect 8162 2694 8176 2746
rect 8200 2694 8214 2746
rect 8214 2694 8226 2746
rect 8226 2694 8256 2746
rect 8280 2694 8290 2746
rect 8290 2694 8336 2746
rect 8040 2692 8096 2694
rect 8120 2692 8176 2694
rect 8200 2692 8256 2694
rect 8280 2692 8336 2694
rect 2628 2202 2684 2204
rect 2708 2202 2764 2204
rect 2788 2202 2844 2204
rect 2868 2202 2924 2204
rect 2628 2150 2674 2202
rect 2674 2150 2684 2202
rect 2708 2150 2738 2202
rect 2738 2150 2750 2202
rect 2750 2150 2764 2202
rect 2788 2150 2802 2202
rect 2802 2150 2814 2202
rect 2814 2150 2844 2202
rect 2868 2150 2878 2202
rect 2878 2150 2924 2202
rect 2628 2148 2684 2150
rect 2708 2148 2764 2150
rect 2788 2148 2844 2150
rect 2868 2148 2924 2150
rect 4652 2202 4708 2204
rect 4732 2202 4788 2204
rect 4812 2202 4868 2204
rect 4892 2202 4948 2204
rect 4652 2150 4698 2202
rect 4698 2150 4708 2202
rect 4732 2150 4762 2202
rect 4762 2150 4774 2202
rect 4774 2150 4788 2202
rect 4812 2150 4826 2202
rect 4826 2150 4838 2202
rect 4838 2150 4868 2202
rect 4892 2150 4902 2202
rect 4902 2150 4948 2202
rect 4652 2148 4708 2150
rect 4732 2148 4788 2150
rect 4812 2148 4868 2150
rect 4892 2148 4948 2150
rect 6676 2202 6732 2204
rect 6756 2202 6812 2204
rect 6836 2202 6892 2204
rect 6916 2202 6972 2204
rect 6676 2150 6722 2202
rect 6722 2150 6732 2202
rect 6756 2150 6786 2202
rect 6786 2150 6798 2202
rect 6798 2150 6812 2202
rect 6836 2150 6850 2202
rect 6850 2150 6862 2202
rect 6862 2150 6892 2202
rect 6916 2150 6926 2202
rect 6926 2150 6972 2202
rect 6676 2148 6732 2150
rect 6756 2148 6812 2150
rect 6836 2148 6892 2150
rect 6916 2148 6972 2150
rect 8700 2202 8756 2204
rect 8780 2202 8836 2204
rect 8860 2202 8916 2204
rect 8940 2202 8996 2204
rect 8700 2150 8746 2202
rect 8746 2150 8756 2202
rect 8780 2150 8810 2202
rect 8810 2150 8822 2202
rect 8822 2150 8836 2202
rect 8860 2150 8874 2202
rect 8874 2150 8886 2202
rect 8886 2150 8916 2202
rect 8940 2150 8950 2202
rect 8950 2150 8996 2202
rect 8700 2148 8756 2150
rect 8780 2148 8836 2150
rect 8860 2148 8916 2150
rect 8940 2148 8996 2150
<< metal3 >>
rect 2618 9824 2934 9825
rect 2618 9760 2624 9824
rect 2688 9760 2704 9824
rect 2768 9760 2784 9824
rect 2848 9760 2864 9824
rect 2928 9760 2934 9824
rect 2618 9759 2934 9760
rect 4642 9824 4958 9825
rect 4642 9760 4648 9824
rect 4712 9760 4728 9824
rect 4792 9760 4808 9824
rect 4872 9760 4888 9824
rect 4952 9760 4958 9824
rect 4642 9759 4958 9760
rect 6666 9824 6982 9825
rect 6666 9760 6672 9824
rect 6736 9760 6752 9824
rect 6816 9760 6832 9824
rect 6896 9760 6912 9824
rect 6976 9760 6982 9824
rect 6666 9759 6982 9760
rect 8690 9824 9006 9825
rect 8690 9760 8696 9824
rect 8760 9760 8776 9824
rect 8840 9760 8856 9824
rect 8920 9760 8936 9824
rect 9000 9760 9006 9824
rect 8690 9759 9006 9760
rect 1958 9280 2274 9281
rect 1958 9216 1964 9280
rect 2028 9216 2044 9280
rect 2108 9216 2124 9280
rect 2188 9216 2204 9280
rect 2268 9216 2274 9280
rect 1958 9215 2274 9216
rect 3982 9280 4298 9281
rect 3982 9216 3988 9280
rect 4052 9216 4068 9280
rect 4132 9216 4148 9280
rect 4212 9216 4228 9280
rect 4292 9216 4298 9280
rect 3982 9215 4298 9216
rect 6006 9280 6322 9281
rect 6006 9216 6012 9280
rect 6076 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6322 9280
rect 6006 9215 6322 9216
rect 8030 9280 8346 9281
rect 8030 9216 8036 9280
rect 8100 9216 8116 9280
rect 8180 9216 8196 9280
rect 8260 9216 8276 9280
rect 8340 9216 8346 9280
rect 8030 9215 8346 9216
rect 0 8938 800 8968
rect 3785 8938 3851 8941
rect 0 8936 3851 8938
rect 0 8880 3790 8936
rect 3846 8880 3851 8936
rect 0 8878 3851 8880
rect 0 8848 800 8878
rect 3785 8875 3851 8878
rect 8661 8938 8727 8941
rect 9517 8938 10317 8968
rect 8661 8936 10317 8938
rect 8661 8880 8666 8936
rect 8722 8880 10317 8936
rect 8661 8878 10317 8880
rect 8661 8875 8727 8878
rect 9517 8848 10317 8878
rect 2618 8736 2934 8737
rect 2618 8672 2624 8736
rect 2688 8672 2704 8736
rect 2768 8672 2784 8736
rect 2848 8672 2864 8736
rect 2928 8672 2934 8736
rect 2618 8671 2934 8672
rect 4642 8736 4958 8737
rect 4642 8672 4648 8736
rect 4712 8672 4728 8736
rect 4792 8672 4808 8736
rect 4872 8672 4888 8736
rect 4952 8672 4958 8736
rect 4642 8671 4958 8672
rect 6666 8736 6982 8737
rect 6666 8672 6672 8736
rect 6736 8672 6752 8736
rect 6816 8672 6832 8736
rect 6896 8672 6912 8736
rect 6976 8672 6982 8736
rect 6666 8671 6982 8672
rect 8690 8736 9006 8737
rect 8690 8672 8696 8736
rect 8760 8672 8776 8736
rect 8840 8672 8856 8736
rect 8920 8672 8936 8736
rect 9000 8672 9006 8736
rect 8690 8671 9006 8672
rect 1958 8192 2274 8193
rect 1958 8128 1964 8192
rect 2028 8128 2044 8192
rect 2108 8128 2124 8192
rect 2188 8128 2204 8192
rect 2268 8128 2274 8192
rect 1958 8127 2274 8128
rect 3982 8192 4298 8193
rect 3982 8128 3988 8192
rect 4052 8128 4068 8192
rect 4132 8128 4148 8192
rect 4212 8128 4228 8192
rect 4292 8128 4298 8192
rect 3982 8127 4298 8128
rect 6006 8192 6322 8193
rect 6006 8128 6012 8192
rect 6076 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6322 8192
rect 6006 8127 6322 8128
rect 8030 8192 8346 8193
rect 8030 8128 8036 8192
rect 8100 8128 8116 8192
rect 8180 8128 8196 8192
rect 8260 8128 8276 8192
rect 8340 8128 8346 8192
rect 8030 8127 8346 8128
rect 3509 7850 3575 7853
rect 4429 7850 4495 7853
rect 3509 7848 4495 7850
rect 3509 7792 3514 7848
rect 3570 7792 4434 7848
rect 4490 7792 4495 7848
rect 3509 7790 4495 7792
rect 3509 7787 3575 7790
rect 4429 7787 4495 7790
rect 2618 7648 2934 7649
rect 0 7578 800 7608
rect 2618 7584 2624 7648
rect 2688 7584 2704 7648
rect 2768 7584 2784 7648
rect 2848 7584 2864 7648
rect 2928 7584 2934 7648
rect 2618 7583 2934 7584
rect 4642 7648 4958 7649
rect 4642 7584 4648 7648
rect 4712 7584 4728 7648
rect 4792 7584 4808 7648
rect 4872 7584 4888 7648
rect 4952 7584 4958 7648
rect 4642 7583 4958 7584
rect 6666 7648 6982 7649
rect 6666 7584 6672 7648
rect 6736 7584 6752 7648
rect 6816 7584 6832 7648
rect 6896 7584 6912 7648
rect 6976 7584 6982 7648
rect 6666 7583 6982 7584
rect 8690 7648 9006 7649
rect 8690 7584 8696 7648
rect 8760 7584 8776 7648
rect 8840 7584 8856 7648
rect 8920 7584 8936 7648
rect 9000 7584 9006 7648
rect 8690 7583 9006 7584
rect 1393 7578 1459 7581
rect 0 7576 1459 7578
rect 0 7520 1398 7576
rect 1454 7520 1459 7576
rect 0 7518 1459 7520
rect 0 7488 800 7518
rect 1393 7515 1459 7518
rect 9121 7578 9187 7581
rect 9517 7578 10317 7608
rect 9121 7576 10317 7578
rect 9121 7520 9126 7576
rect 9182 7520 10317 7576
rect 9121 7518 10317 7520
rect 9121 7515 9187 7518
rect 9517 7488 10317 7518
rect 1958 7104 2274 7105
rect 1958 7040 1964 7104
rect 2028 7040 2044 7104
rect 2108 7040 2124 7104
rect 2188 7040 2204 7104
rect 2268 7040 2274 7104
rect 1958 7039 2274 7040
rect 3982 7104 4298 7105
rect 3982 7040 3988 7104
rect 4052 7040 4068 7104
rect 4132 7040 4148 7104
rect 4212 7040 4228 7104
rect 4292 7040 4298 7104
rect 3982 7039 4298 7040
rect 6006 7104 6322 7105
rect 6006 7040 6012 7104
rect 6076 7040 6092 7104
rect 6156 7040 6172 7104
rect 6236 7040 6252 7104
rect 6316 7040 6322 7104
rect 6006 7039 6322 7040
rect 8030 7104 8346 7105
rect 8030 7040 8036 7104
rect 8100 7040 8116 7104
rect 8180 7040 8196 7104
rect 8260 7040 8276 7104
rect 8340 7040 8346 7104
rect 8030 7039 8346 7040
rect 8569 6898 8635 6901
rect 9517 6898 10317 6928
rect 8569 6896 10317 6898
rect 8569 6840 8574 6896
rect 8630 6840 10317 6896
rect 8569 6838 10317 6840
rect 8569 6835 8635 6838
rect 9517 6808 10317 6838
rect 2618 6560 2934 6561
rect 2618 6496 2624 6560
rect 2688 6496 2704 6560
rect 2768 6496 2784 6560
rect 2848 6496 2864 6560
rect 2928 6496 2934 6560
rect 2618 6495 2934 6496
rect 4642 6560 4958 6561
rect 4642 6496 4648 6560
rect 4712 6496 4728 6560
rect 4792 6496 4808 6560
rect 4872 6496 4888 6560
rect 4952 6496 4958 6560
rect 4642 6495 4958 6496
rect 6666 6560 6982 6561
rect 6666 6496 6672 6560
rect 6736 6496 6752 6560
rect 6816 6496 6832 6560
rect 6896 6496 6912 6560
rect 6976 6496 6982 6560
rect 6666 6495 6982 6496
rect 8690 6560 9006 6561
rect 8690 6496 8696 6560
rect 8760 6496 8776 6560
rect 8840 6496 8856 6560
rect 8920 6496 8936 6560
rect 9000 6496 9006 6560
rect 8690 6495 9006 6496
rect 0 6218 800 6248
rect 8661 6218 8727 6221
rect 9517 6218 10317 6248
rect 0 6128 858 6218
rect 8661 6216 10317 6218
rect 8661 6160 8666 6216
rect 8722 6160 10317 6216
rect 8661 6158 10317 6160
rect 8661 6155 8727 6158
rect 9517 6128 10317 6158
rect 798 5949 858 6128
rect 1958 6016 2274 6017
rect 1958 5952 1964 6016
rect 2028 5952 2044 6016
rect 2108 5952 2124 6016
rect 2188 5952 2204 6016
rect 2268 5952 2274 6016
rect 1958 5951 2274 5952
rect 3982 6016 4298 6017
rect 3982 5952 3988 6016
rect 4052 5952 4068 6016
rect 4132 5952 4148 6016
rect 4212 5952 4228 6016
rect 4292 5952 4298 6016
rect 3982 5951 4298 5952
rect 6006 6016 6322 6017
rect 6006 5952 6012 6016
rect 6076 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6322 6016
rect 6006 5951 6322 5952
rect 8030 6016 8346 6017
rect 8030 5952 8036 6016
rect 8100 5952 8116 6016
rect 8180 5952 8196 6016
rect 8260 5952 8276 6016
rect 8340 5952 8346 6016
rect 8030 5951 8346 5952
rect 749 5944 858 5949
rect 749 5888 754 5944
rect 810 5888 858 5944
rect 749 5886 858 5888
rect 749 5883 815 5886
rect 2618 5472 2934 5473
rect 2618 5408 2624 5472
rect 2688 5408 2704 5472
rect 2768 5408 2784 5472
rect 2848 5408 2864 5472
rect 2928 5408 2934 5472
rect 2618 5407 2934 5408
rect 4642 5472 4958 5473
rect 4642 5408 4648 5472
rect 4712 5408 4728 5472
rect 4792 5408 4808 5472
rect 4872 5408 4888 5472
rect 4952 5408 4958 5472
rect 4642 5407 4958 5408
rect 6666 5472 6982 5473
rect 6666 5408 6672 5472
rect 6736 5408 6752 5472
rect 6816 5408 6832 5472
rect 6896 5408 6912 5472
rect 6976 5408 6982 5472
rect 6666 5407 6982 5408
rect 8690 5472 9006 5473
rect 8690 5408 8696 5472
rect 8760 5408 8776 5472
rect 8840 5408 8856 5472
rect 8920 5408 8936 5472
rect 9000 5408 9006 5472
rect 8690 5407 9006 5408
rect 1958 4928 2274 4929
rect 1958 4864 1964 4928
rect 2028 4864 2044 4928
rect 2108 4864 2124 4928
rect 2188 4864 2204 4928
rect 2268 4864 2274 4928
rect 1958 4863 2274 4864
rect 3982 4928 4298 4929
rect 3982 4864 3988 4928
rect 4052 4864 4068 4928
rect 4132 4864 4148 4928
rect 4212 4864 4228 4928
rect 4292 4864 4298 4928
rect 3982 4863 4298 4864
rect 6006 4928 6322 4929
rect 6006 4864 6012 4928
rect 6076 4864 6092 4928
rect 6156 4864 6172 4928
rect 6236 4864 6252 4928
rect 6316 4864 6322 4928
rect 6006 4863 6322 4864
rect 8030 4928 8346 4929
rect 8030 4864 8036 4928
rect 8100 4864 8116 4928
rect 8180 4864 8196 4928
rect 8260 4864 8276 4928
rect 8340 4864 8346 4928
rect 8030 4863 8346 4864
rect 8753 4858 8819 4861
rect 9517 4858 10317 4888
rect 8753 4856 10317 4858
rect 8753 4800 8758 4856
rect 8814 4800 10317 4856
rect 8753 4798 10317 4800
rect 8753 4795 8819 4798
rect 9517 4768 10317 4798
rect 2618 4384 2934 4385
rect 2618 4320 2624 4384
rect 2688 4320 2704 4384
rect 2768 4320 2784 4384
rect 2848 4320 2864 4384
rect 2928 4320 2934 4384
rect 2618 4319 2934 4320
rect 4642 4384 4958 4385
rect 4642 4320 4648 4384
rect 4712 4320 4728 4384
rect 4792 4320 4808 4384
rect 4872 4320 4888 4384
rect 4952 4320 4958 4384
rect 4642 4319 4958 4320
rect 6666 4384 6982 4385
rect 6666 4320 6672 4384
rect 6736 4320 6752 4384
rect 6816 4320 6832 4384
rect 6896 4320 6912 4384
rect 6976 4320 6982 4384
rect 6666 4319 6982 4320
rect 8690 4384 9006 4385
rect 8690 4320 8696 4384
rect 8760 4320 8776 4384
rect 8840 4320 8856 4384
rect 8920 4320 8936 4384
rect 9000 4320 9006 4384
rect 8690 4319 9006 4320
rect 9121 4178 9187 4181
rect 9517 4178 10317 4208
rect 9121 4176 10317 4178
rect 9121 4120 9126 4176
rect 9182 4120 10317 4176
rect 9121 4118 10317 4120
rect 9121 4115 9187 4118
rect 9517 4088 10317 4118
rect 1958 3840 2274 3841
rect 1958 3776 1964 3840
rect 2028 3776 2044 3840
rect 2108 3776 2124 3840
rect 2188 3776 2204 3840
rect 2268 3776 2274 3840
rect 1958 3775 2274 3776
rect 3982 3840 4298 3841
rect 3982 3776 3988 3840
rect 4052 3776 4068 3840
rect 4132 3776 4148 3840
rect 4212 3776 4228 3840
rect 4292 3776 4298 3840
rect 3982 3775 4298 3776
rect 6006 3840 6322 3841
rect 6006 3776 6012 3840
rect 6076 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6322 3840
rect 6006 3775 6322 3776
rect 8030 3840 8346 3841
rect 8030 3776 8036 3840
rect 8100 3776 8116 3840
rect 8180 3776 8196 3840
rect 8260 3776 8276 3840
rect 8340 3776 8346 3840
rect 8030 3775 8346 3776
rect 8661 3498 8727 3501
rect 9517 3498 10317 3528
rect 8661 3496 10317 3498
rect 8661 3440 8666 3496
rect 8722 3440 10317 3496
rect 8661 3438 10317 3440
rect 8661 3435 8727 3438
rect 9517 3408 10317 3438
rect 2618 3296 2934 3297
rect 2618 3232 2624 3296
rect 2688 3232 2704 3296
rect 2768 3232 2784 3296
rect 2848 3232 2864 3296
rect 2928 3232 2934 3296
rect 2618 3231 2934 3232
rect 4642 3296 4958 3297
rect 4642 3232 4648 3296
rect 4712 3232 4728 3296
rect 4792 3232 4808 3296
rect 4872 3232 4888 3296
rect 4952 3232 4958 3296
rect 4642 3231 4958 3232
rect 6666 3296 6982 3297
rect 6666 3232 6672 3296
rect 6736 3232 6752 3296
rect 6816 3232 6832 3296
rect 6896 3232 6912 3296
rect 6976 3232 6982 3296
rect 6666 3231 6982 3232
rect 8690 3296 9006 3297
rect 8690 3232 8696 3296
rect 8760 3232 8776 3296
rect 8840 3232 8856 3296
rect 8920 3232 8936 3296
rect 9000 3232 9006 3296
rect 8690 3231 9006 3232
rect 8753 2818 8819 2821
rect 9517 2818 10317 2848
rect 8753 2816 10317 2818
rect 8753 2760 8758 2816
rect 8814 2760 10317 2816
rect 8753 2758 10317 2760
rect 8753 2755 8819 2758
rect 1958 2752 2274 2753
rect 1958 2688 1964 2752
rect 2028 2688 2044 2752
rect 2108 2688 2124 2752
rect 2188 2688 2204 2752
rect 2268 2688 2274 2752
rect 1958 2687 2274 2688
rect 3982 2752 4298 2753
rect 3982 2688 3988 2752
rect 4052 2688 4068 2752
rect 4132 2688 4148 2752
rect 4212 2688 4228 2752
rect 4292 2688 4298 2752
rect 3982 2687 4298 2688
rect 6006 2752 6322 2753
rect 6006 2688 6012 2752
rect 6076 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6322 2752
rect 6006 2687 6322 2688
rect 8030 2752 8346 2753
rect 8030 2688 8036 2752
rect 8100 2688 8116 2752
rect 8180 2688 8196 2752
rect 8260 2688 8276 2752
rect 8340 2688 8346 2752
rect 9517 2728 10317 2758
rect 8030 2687 8346 2688
rect 2618 2208 2934 2209
rect 2618 2144 2624 2208
rect 2688 2144 2704 2208
rect 2768 2144 2784 2208
rect 2848 2144 2864 2208
rect 2928 2144 2934 2208
rect 2618 2143 2934 2144
rect 4642 2208 4958 2209
rect 4642 2144 4648 2208
rect 4712 2144 4728 2208
rect 4792 2144 4808 2208
rect 4872 2144 4888 2208
rect 4952 2144 4958 2208
rect 4642 2143 4958 2144
rect 6666 2208 6982 2209
rect 6666 2144 6672 2208
rect 6736 2144 6752 2208
rect 6816 2144 6832 2208
rect 6896 2144 6912 2208
rect 6976 2144 6982 2208
rect 6666 2143 6982 2144
rect 8690 2208 9006 2209
rect 8690 2144 8696 2208
rect 8760 2144 8776 2208
rect 8840 2144 8856 2208
rect 8920 2144 8936 2208
rect 9000 2144 9006 2208
rect 8690 2143 9006 2144
<< via3 >>
rect 2624 9820 2688 9824
rect 2624 9764 2628 9820
rect 2628 9764 2684 9820
rect 2684 9764 2688 9820
rect 2624 9760 2688 9764
rect 2704 9820 2768 9824
rect 2704 9764 2708 9820
rect 2708 9764 2764 9820
rect 2764 9764 2768 9820
rect 2704 9760 2768 9764
rect 2784 9820 2848 9824
rect 2784 9764 2788 9820
rect 2788 9764 2844 9820
rect 2844 9764 2848 9820
rect 2784 9760 2848 9764
rect 2864 9820 2928 9824
rect 2864 9764 2868 9820
rect 2868 9764 2924 9820
rect 2924 9764 2928 9820
rect 2864 9760 2928 9764
rect 4648 9820 4712 9824
rect 4648 9764 4652 9820
rect 4652 9764 4708 9820
rect 4708 9764 4712 9820
rect 4648 9760 4712 9764
rect 4728 9820 4792 9824
rect 4728 9764 4732 9820
rect 4732 9764 4788 9820
rect 4788 9764 4792 9820
rect 4728 9760 4792 9764
rect 4808 9820 4872 9824
rect 4808 9764 4812 9820
rect 4812 9764 4868 9820
rect 4868 9764 4872 9820
rect 4808 9760 4872 9764
rect 4888 9820 4952 9824
rect 4888 9764 4892 9820
rect 4892 9764 4948 9820
rect 4948 9764 4952 9820
rect 4888 9760 4952 9764
rect 6672 9820 6736 9824
rect 6672 9764 6676 9820
rect 6676 9764 6732 9820
rect 6732 9764 6736 9820
rect 6672 9760 6736 9764
rect 6752 9820 6816 9824
rect 6752 9764 6756 9820
rect 6756 9764 6812 9820
rect 6812 9764 6816 9820
rect 6752 9760 6816 9764
rect 6832 9820 6896 9824
rect 6832 9764 6836 9820
rect 6836 9764 6892 9820
rect 6892 9764 6896 9820
rect 6832 9760 6896 9764
rect 6912 9820 6976 9824
rect 6912 9764 6916 9820
rect 6916 9764 6972 9820
rect 6972 9764 6976 9820
rect 6912 9760 6976 9764
rect 8696 9820 8760 9824
rect 8696 9764 8700 9820
rect 8700 9764 8756 9820
rect 8756 9764 8760 9820
rect 8696 9760 8760 9764
rect 8776 9820 8840 9824
rect 8776 9764 8780 9820
rect 8780 9764 8836 9820
rect 8836 9764 8840 9820
rect 8776 9760 8840 9764
rect 8856 9820 8920 9824
rect 8856 9764 8860 9820
rect 8860 9764 8916 9820
rect 8916 9764 8920 9820
rect 8856 9760 8920 9764
rect 8936 9820 9000 9824
rect 8936 9764 8940 9820
rect 8940 9764 8996 9820
rect 8996 9764 9000 9820
rect 8936 9760 9000 9764
rect 1964 9276 2028 9280
rect 1964 9220 1968 9276
rect 1968 9220 2024 9276
rect 2024 9220 2028 9276
rect 1964 9216 2028 9220
rect 2044 9276 2108 9280
rect 2044 9220 2048 9276
rect 2048 9220 2104 9276
rect 2104 9220 2108 9276
rect 2044 9216 2108 9220
rect 2124 9276 2188 9280
rect 2124 9220 2128 9276
rect 2128 9220 2184 9276
rect 2184 9220 2188 9276
rect 2124 9216 2188 9220
rect 2204 9276 2268 9280
rect 2204 9220 2208 9276
rect 2208 9220 2264 9276
rect 2264 9220 2268 9276
rect 2204 9216 2268 9220
rect 3988 9276 4052 9280
rect 3988 9220 3992 9276
rect 3992 9220 4048 9276
rect 4048 9220 4052 9276
rect 3988 9216 4052 9220
rect 4068 9276 4132 9280
rect 4068 9220 4072 9276
rect 4072 9220 4128 9276
rect 4128 9220 4132 9276
rect 4068 9216 4132 9220
rect 4148 9276 4212 9280
rect 4148 9220 4152 9276
rect 4152 9220 4208 9276
rect 4208 9220 4212 9276
rect 4148 9216 4212 9220
rect 4228 9276 4292 9280
rect 4228 9220 4232 9276
rect 4232 9220 4288 9276
rect 4288 9220 4292 9276
rect 4228 9216 4292 9220
rect 6012 9276 6076 9280
rect 6012 9220 6016 9276
rect 6016 9220 6072 9276
rect 6072 9220 6076 9276
rect 6012 9216 6076 9220
rect 6092 9276 6156 9280
rect 6092 9220 6096 9276
rect 6096 9220 6152 9276
rect 6152 9220 6156 9276
rect 6092 9216 6156 9220
rect 6172 9276 6236 9280
rect 6172 9220 6176 9276
rect 6176 9220 6232 9276
rect 6232 9220 6236 9276
rect 6172 9216 6236 9220
rect 6252 9276 6316 9280
rect 6252 9220 6256 9276
rect 6256 9220 6312 9276
rect 6312 9220 6316 9276
rect 6252 9216 6316 9220
rect 8036 9276 8100 9280
rect 8036 9220 8040 9276
rect 8040 9220 8096 9276
rect 8096 9220 8100 9276
rect 8036 9216 8100 9220
rect 8116 9276 8180 9280
rect 8116 9220 8120 9276
rect 8120 9220 8176 9276
rect 8176 9220 8180 9276
rect 8116 9216 8180 9220
rect 8196 9276 8260 9280
rect 8196 9220 8200 9276
rect 8200 9220 8256 9276
rect 8256 9220 8260 9276
rect 8196 9216 8260 9220
rect 8276 9276 8340 9280
rect 8276 9220 8280 9276
rect 8280 9220 8336 9276
rect 8336 9220 8340 9276
rect 8276 9216 8340 9220
rect 2624 8732 2688 8736
rect 2624 8676 2628 8732
rect 2628 8676 2684 8732
rect 2684 8676 2688 8732
rect 2624 8672 2688 8676
rect 2704 8732 2768 8736
rect 2704 8676 2708 8732
rect 2708 8676 2764 8732
rect 2764 8676 2768 8732
rect 2704 8672 2768 8676
rect 2784 8732 2848 8736
rect 2784 8676 2788 8732
rect 2788 8676 2844 8732
rect 2844 8676 2848 8732
rect 2784 8672 2848 8676
rect 2864 8732 2928 8736
rect 2864 8676 2868 8732
rect 2868 8676 2924 8732
rect 2924 8676 2928 8732
rect 2864 8672 2928 8676
rect 4648 8732 4712 8736
rect 4648 8676 4652 8732
rect 4652 8676 4708 8732
rect 4708 8676 4712 8732
rect 4648 8672 4712 8676
rect 4728 8732 4792 8736
rect 4728 8676 4732 8732
rect 4732 8676 4788 8732
rect 4788 8676 4792 8732
rect 4728 8672 4792 8676
rect 4808 8732 4872 8736
rect 4808 8676 4812 8732
rect 4812 8676 4868 8732
rect 4868 8676 4872 8732
rect 4808 8672 4872 8676
rect 4888 8732 4952 8736
rect 4888 8676 4892 8732
rect 4892 8676 4948 8732
rect 4948 8676 4952 8732
rect 4888 8672 4952 8676
rect 6672 8732 6736 8736
rect 6672 8676 6676 8732
rect 6676 8676 6732 8732
rect 6732 8676 6736 8732
rect 6672 8672 6736 8676
rect 6752 8732 6816 8736
rect 6752 8676 6756 8732
rect 6756 8676 6812 8732
rect 6812 8676 6816 8732
rect 6752 8672 6816 8676
rect 6832 8732 6896 8736
rect 6832 8676 6836 8732
rect 6836 8676 6892 8732
rect 6892 8676 6896 8732
rect 6832 8672 6896 8676
rect 6912 8732 6976 8736
rect 6912 8676 6916 8732
rect 6916 8676 6972 8732
rect 6972 8676 6976 8732
rect 6912 8672 6976 8676
rect 8696 8732 8760 8736
rect 8696 8676 8700 8732
rect 8700 8676 8756 8732
rect 8756 8676 8760 8732
rect 8696 8672 8760 8676
rect 8776 8732 8840 8736
rect 8776 8676 8780 8732
rect 8780 8676 8836 8732
rect 8836 8676 8840 8732
rect 8776 8672 8840 8676
rect 8856 8732 8920 8736
rect 8856 8676 8860 8732
rect 8860 8676 8916 8732
rect 8916 8676 8920 8732
rect 8856 8672 8920 8676
rect 8936 8732 9000 8736
rect 8936 8676 8940 8732
rect 8940 8676 8996 8732
rect 8996 8676 9000 8732
rect 8936 8672 9000 8676
rect 1964 8188 2028 8192
rect 1964 8132 1968 8188
rect 1968 8132 2024 8188
rect 2024 8132 2028 8188
rect 1964 8128 2028 8132
rect 2044 8188 2108 8192
rect 2044 8132 2048 8188
rect 2048 8132 2104 8188
rect 2104 8132 2108 8188
rect 2044 8128 2108 8132
rect 2124 8188 2188 8192
rect 2124 8132 2128 8188
rect 2128 8132 2184 8188
rect 2184 8132 2188 8188
rect 2124 8128 2188 8132
rect 2204 8188 2268 8192
rect 2204 8132 2208 8188
rect 2208 8132 2264 8188
rect 2264 8132 2268 8188
rect 2204 8128 2268 8132
rect 3988 8188 4052 8192
rect 3988 8132 3992 8188
rect 3992 8132 4048 8188
rect 4048 8132 4052 8188
rect 3988 8128 4052 8132
rect 4068 8188 4132 8192
rect 4068 8132 4072 8188
rect 4072 8132 4128 8188
rect 4128 8132 4132 8188
rect 4068 8128 4132 8132
rect 4148 8188 4212 8192
rect 4148 8132 4152 8188
rect 4152 8132 4208 8188
rect 4208 8132 4212 8188
rect 4148 8128 4212 8132
rect 4228 8188 4292 8192
rect 4228 8132 4232 8188
rect 4232 8132 4288 8188
rect 4288 8132 4292 8188
rect 4228 8128 4292 8132
rect 6012 8188 6076 8192
rect 6012 8132 6016 8188
rect 6016 8132 6072 8188
rect 6072 8132 6076 8188
rect 6012 8128 6076 8132
rect 6092 8188 6156 8192
rect 6092 8132 6096 8188
rect 6096 8132 6152 8188
rect 6152 8132 6156 8188
rect 6092 8128 6156 8132
rect 6172 8188 6236 8192
rect 6172 8132 6176 8188
rect 6176 8132 6232 8188
rect 6232 8132 6236 8188
rect 6172 8128 6236 8132
rect 6252 8188 6316 8192
rect 6252 8132 6256 8188
rect 6256 8132 6312 8188
rect 6312 8132 6316 8188
rect 6252 8128 6316 8132
rect 8036 8188 8100 8192
rect 8036 8132 8040 8188
rect 8040 8132 8096 8188
rect 8096 8132 8100 8188
rect 8036 8128 8100 8132
rect 8116 8188 8180 8192
rect 8116 8132 8120 8188
rect 8120 8132 8176 8188
rect 8176 8132 8180 8188
rect 8116 8128 8180 8132
rect 8196 8188 8260 8192
rect 8196 8132 8200 8188
rect 8200 8132 8256 8188
rect 8256 8132 8260 8188
rect 8196 8128 8260 8132
rect 8276 8188 8340 8192
rect 8276 8132 8280 8188
rect 8280 8132 8336 8188
rect 8336 8132 8340 8188
rect 8276 8128 8340 8132
rect 2624 7644 2688 7648
rect 2624 7588 2628 7644
rect 2628 7588 2684 7644
rect 2684 7588 2688 7644
rect 2624 7584 2688 7588
rect 2704 7644 2768 7648
rect 2704 7588 2708 7644
rect 2708 7588 2764 7644
rect 2764 7588 2768 7644
rect 2704 7584 2768 7588
rect 2784 7644 2848 7648
rect 2784 7588 2788 7644
rect 2788 7588 2844 7644
rect 2844 7588 2848 7644
rect 2784 7584 2848 7588
rect 2864 7644 2928 7648
rect 2864 7588 2868 7644
rect 2868 7588 2924 7644
rect 2924 7588 2928 7644
rect 2864 7584 2928 7588
rect 4648 7644 4712 7648
rect 4648 7588 4652 7644
rect 4652 7588 4708 7644
rect 4708 7588 4712 7644
rect 4648 7584 4712 7588
rect 4728 7644 4792 7648
rect 4728 7588 4732 7644
rect 4732 7588 4788 7644
rect 4788 7588 4792 7644
rect 4728 7584 4792 7588
rect 4808 7644 4872 7648
rect 4808 7588 4812 7644
rect 4812 7588 4868 7644
rect 4868 7588 4872 7644
rect 4808 7584 4872 7588
rect 4888 7644 4952 7648
rect 4888 7588 4892 7644
rect 4892 7588 4948 7644
rect 4948 7588 4952 7644
rect 4888 7584 4952 7588
rect 6672 7644 6736 7648
rect 6672 7588 6676 7644
rect 6676 7588 6732 7644
rect 6732 7588 6736 7644
rect 6672 7584 6736 7588
rect 6752 7644 6816 7648
rect 6752 7588 6756 7644
rect 6756 7588 6812 7644
rect 6812 7588 6816 7644
rect 6752 7584 6816 7588
rect 6832 7644 6896 7648
rect 6832 7588 6836 7644
rect 6836 7588 6892 7644
rect 6892 7588 6896 7644
rect 6832 7584 6896 7588
rect 6912 7644 6976 7648
rect 6912 7588 6916 7644
rect 6916 7588 6972 7644
rect 6972 7588 6976 7644
rect 6912 7584 6976 7588
rect 8696 7644 8760 7648
rect 8696 7588 8700 7644
rect 8700 7588 8756 7644
rect 8756 7588 8760 7644
rect 8696 7584 8760 7588
rect 8776 7644 8840 7648
rect 8776 7588 8780 7644
rect 8780 7588 8836 7644
rect 8836 7588 8840 7644
rect 8776 7584 8840 7588
rect 8856 7644 8920 7648
rect 8856 7588 8860 7644
rect 8860 7588 8916 7644
rect 8916 7588 8920 7644
rect 8856 7584 8920 7588
rect 8936 7644 9000 7648
rect 8936 7588 8940 7644
rect 8940 7588 8996 7644
rect 8996 7588 9000 7644
rect 8936 7584 9000 7588
rect 1964 7100 2028 7104
rect 1964 7044 1968 7100
rect 1968 7044 2024 7100
rect 2024 7044 2028 7100
rect 1964 7040 2028 7044
rect 2044 7100 2108 7104
rect 2044 7044 2048 7100
rect 2048 7044 2104 7100
rect 2104 7044 2108 7100
rect 2044 7040 2108 7044
rect 2124 7100 2188 7104
rect 2124 7044 2128 7100
rect 2128 7044 2184 7100
rect 2184 7044 2188 7100
rect 2124 7040 2188 7044
rect 2204 7100 2268 7104
rect 2204 7044 2208 7100
rect 2208 7044 2264 7100
rect 2264 7044 2268 7100
rect 2204 7040 2268 7044
rect 3988 7100 4052 7104
rect 3988 7044 3992 7100
rect 3992 7044 4048 7100
rect 4048 7044 4052 7100
rect 3988 7040 4052 7044
rect 4068 7100 4132 7104
rect 4068 7044 4072 7100
rect 4072 7044 4128 7100
rect 4128 7044 4132 7100
rect 4068 7040 4132 7044
rect 4148 7100 4212 7104
rect 4148 7044 4152 7100
rect 4152 7044 4208 7100
rect 4208 7044 4212 7100
rect 4148 7040 4212 7044
rect 4228 7100 4292 7104
rect 4228 7044 4232 7100
rect 4232 7044 4288 7100
rect 4288 7044 4292 7100
rect 4228 7040 4292 7044
rect 6012 7100 6076 7104
rect 6012 7044 6016 7100
rect 6016 7044 6072 7100
rect 6072 7044 6076 7100
rect 6012 7040 6076 7044
rect 6092 7100 6156 7104
rect 6092 7044 6096 7100
rect 6096 7044 6152 7100
rect 6152 7044 6156 7100
rect 6092 7040 6156 7044
rect 6172 7100 6236 7104
rect 6172 7044 6176 7100
rect 6176 7044 6232 7100
rect 6232 7044 6236 7100
rect 6172 7040 6236 7044
rect 6252 7100 6316 7104
rect 6252 7044 6256 7100
rect 6256 7044 6312 7100
rect 6312 7044 6316 7100
rect 6252 7040 6316 7044
rect 8036 7100 8100 7104
rect 8036 7044 8040 7100
rect 8040 7044 8096 7100
rect 8096 7044 8100 7100
rect 8036 7040 8100 7044
rect 8116 7100 8180 7104
rect 8116 7044 8120 7100
rect 8120 7044 8176 7100
rect 8176 7044 8180 7100
rect 8116 7040 8180 7044
rect 8196 7100 8260 7104
rect 8196 7044 8200 7100
rect 8200 7044 8256 7100
rect 8256 7044 8260 7100
rect 8196 7040 8260 7044
rect 8276 7100 8340 7104
rect 8276 7044 8280 7100
rect 8280 7044 8336 7100
rect 8336 7044 8340 7100
rect 8276 7040 8340 7044
rect 2624 6556 2688 6560
rect 2624 6500 2628 6556
rect 2628 6500 2684 6556
rect 2684 6500 2688 6556
rect 2624 6496 2688 6500
rect 2704 6556 2768 6560
rect 2704 6500 2708 6556
rect 2708 6500 2764 6556
rect 2764 6500 2768 6556
rect 2704 6496 2768 6500
rect 2784 6556 2848 6560
rect 2784 6500 2788 6556
rect 2788 6500 2844 6556
rect 2844 6500 2848 6556
rect 2784 6496 2848 6500
rect 2864 6556 2928 6560
rect 2864 6500 2868 6556
rect 2868 6500 2924 6556
rect 2924 6500 2928 6556
rect 2864 6496 2928 6500
rect 4648 6556 4712 6560
rect 4648 6500 4652 6556
rect 4652 6500 4708 6556
rect 4708 6500 4712 6556
rect 4648 6496 4712 6500
rect 4728 6556 4792 6560
rect 4728 6500 4732 6556
rect 4732 6500 4788 6556
rect 4788 6500 4792 6556
rect 4728 6496 4792 6500
rect 4808 6556 4872 6560
rect 4808 6500 4812 6556
rect 4812 6500 4868 6556
rect 4868 6500 4872 6556
rect 4808 6496 4872 6500
rect 4888 6556 4952 6560
rect 4888 6500 4892 6556
rect 4892 6500 4948 6556
rect 4948 6500 4952 6556
rect 4888 6496 4952 6500
rect 6672 6556 6736 6560
rect 6672 6500 6676 6556
rect 6676 6500 6732 6556
rect 6732 6500 6736 6556
rect 6672 6496 6736 6500
rect 6752 6556 6816 6560
rect 6752 6500 6756 6556
rect 6756 6500 6812 6556
rect 6812 6500 6816 6556
rect 6752 6496 6816 6500
rect 6832 6556 6896 6560
rect 6832 6500 6836 6556
rect 6836 6500 6892 6556
rect 6892 6500 6896 6556
rect 6832 6496 6896 6500
rect 6912 6556 6976 6560
rect 6912 6500 6916 6556
rect 6916 6500 6972 6556
rect 6972 6500 6976 6556
rect 6912 6496 6976 6500
rect 8696 6556 8760 6560
rect 8696 6500 8700 6556
rect 8700 6500 8756 6556
rect 8756 6500 8760 6556
rect 8696 6496 8760 6500
rect 8776 6556 8840 6560
rect 8776 6500 8780 6556
rect 8780 6500 8836 6556
rect 8836 6500 8840 6556
rect 8776 6496 8840 6500
rect 8856 6556 8920 6560
rect 8856 6500 8860 6556
rect 8860 6500 8916 6556
rect 8916 6500 8920 6556
rect 8856 6496 8920 6500
rect 8936 6556 9000 6560
rect 8936 6500 8940 6556
rect 8940 6500 8996 6556
rect 8996 6500 9000 6556
rect 8936 6496 9000 6500
rect 1964 6012 2028 6016
rect 1964 5956 1968 6012
rect 1968 5956 2024 6012
rect 2024 5956 2028 6012
rect 1964 5952 2028 5956
rect 2044 6012 2108 6016
rect 2044 5956 2048 6012
rect 2048 5956 2104 6012
rect 2104 5956 2108 6012
rect 2044 5952 2108 5956
rect 2124 6012 2188 6016
rect 2124 5956 2128 6012
rect 2128 5956 2184 6012
rect 2184 5956 2188 6012
rect 2124 5952 2188 5956
rect 2204 6012 2268 6016
rect 2204 5956 2208 6012
rect 2208 5956 2264 6012
rect 2264 5956 2268 6012
rect 2204 5952 2268 5956
rect 3988 6012 4052 6016
rect 3988 5956 3992 6012
rect 3992 5956 4048 6012
rect 4048 5956 4052 6012
rect 3988 5952 4052 5956
rect 4068 6012 4132 6016
rect 4068 5956 4072 6012
rect 4072 5956 4128 6012
rect 4128 5956 4132 6012
rect 4068 5952 4132 5956
rect 4148 6012 4212 6016
rect 4148 5956 4152 6012
rect 4152 5956 4208 6012
rect 4208 5956 4212 6012
rect 4148 5952 4212 5956
rect 4228 6012 4292 6016
rect 4228 5956 4232 6012
rect 4232 5956 4288 6012
rect 4288 5956 4292 6012
rect 4228 5952 4292 5956
rect 6012 6012 6076 6016
rect 6012 5956 6016 6012
rect 6016 5956 6072 6012
rect 6072 5956 6076 6012
rect 6012 5952 6076 5956
rect 6092 6012 6156 6016
rect 6092 5956 6096 6012
rect 6096 5956 6152 6012
rect 6152 5956 6156 6012
rect 6092 5952 6156 5956
rect 6172 6012 6236 6016
rect 6172 5956 6176 6012
rect 6176 5956 6232 6012
rect 6232 5956 6236 6012
rect 6172 5952 6236 5956
rect 6252 6012 6316 6016
rect 6252 5956 6256 6012
rect 6256 5956 6312 6012
rect 6312 5956 6316 6012
rect 6252 5952 6316 5956
rect 8036 6012 8100 6016
rect 8036 5956 8040 6012
rect 8040 5956 8096 6012
rect 8096 5956 8100 6012
rect 8036 5952 8100 5956
rect 8116 6012 8180 6016
rect 8116 5956 8120 6012
rect 8120 5956 8176 6012
rect 8176 5956 8180 6012
rect 8116 5952 8180 5956
rect 8196 6012 8260 6016
rect 8196 5956 8200 6012
rect 8200 5956 8256 6012
rect 8256 5956 8260 6012
rect 8196 5952 8260 5956
rect 8276 6012 8340 6016
rect 8276 5956 8280 6012
rect 8280 5956 8336 6012
rect 8336 5956 8340 6012
rect 8276 5952 8340 5956
rect 2624 5468 2688 5472
rect 2624 5412 2628 5468
rect 2628 5412 2684 5468
rect 2684 5412 2688 5468
rect 2624 5408 2688 5412
rect 2704 5468 2768 5472
rect 2704 5412 2708 5468
rect 2708 5412 2764 5468
rect 2764 5412 2768 5468
rect 2704 5408 2768 5412
rect 2784 5468 2848 5472
rect 2784 5412 2788 5468
rect 2788 5412 2844 5468
rect 2844 5412 2848 5468
rect 2784 5408 2848 5412
rect 2864 5468 2928 5472
rect 2864 5412 2868 5468
rect 2868 5412 2924 5468
rect 2924 5412 2928 5468
rect 2864 5408 2928 5412
rect 4648 5468 4712 5472
rect 4648 5412 4652 5468
rect 4652 5412 4708 5468
rect 4708 5412 4712 5468
rect 4648 5408 4712 5412
rect 4728 5468 4792 5472
rect 4728 5412 4732 5468
rect 4732 5412 4788 5468
rect 4788 5412 4792 5468
rect 4728 5408 4792 5412
rect 4808 5468 4872 5472
rect 4808 5412 4812 5468
rect 4812 5412 4868 5468
rect 4868 5412 4872 5468
rect 4808 5408 4872 5412
rect 4888 5468 4952 5472
rect 4888 5412 4892 5468
rect 4892 5412 4948 5468
rect 4948 5412 4952 5468
rect 4888 5408 4952 5412
rect 6672 5468 6736 5472
rect 6672 5412 6676 5468
rect 6676 5412 6732 5468
rect 6732 5412 6736 5468
rect 6672 5408 6736 5412
rect 6752 5468 6816 5472
rect 6752 5412 6756 5468
rect 6756 5412 6812 5468
rect 6812 5412 6816 5468
rect 6752 5408 6816 5412
rect 6832 5468 6896 5472
rect 6832 5412 6836 5468
rect 6836 5412 6892 5468
rect 6892 5412 6896 5468
rect 6832 5408 6896 5412
rect 6912 5468 6976 5472
rect 6912 5412 6916 5468
rect 6916 5412 6972 5468
rect 6972 5412 6976 5468
rect 6912 5408 6976 5412
rect 8696 5468 8760 5472
rect 8696 5412 8700 5468
rect 8700 5412 8756 5468
rect 8756 5412 8760 5468
rect 8696 5408 8760 5412
rect 8776 5468 8840 5472
rect 8776 5412 8780 5468
rect 8780 5412 8836 5468
rect 8836 5412 8840 5468
rect 8776 5408 8840 5412
rect 8856 5468 8920 5472
rect 8856 5412 8860 5468
rect 8860 5412 8916 5468
rect 8916 5412 8920 5468
rect 8856 5408 8920 5412
rect 8936 5468 9000 5472
rect 8936 5412 8940 5468
rect 8940 5412 8996 5468
rect 8996 5412 9000 5468
rect 8936 5408 9000 5412
rect 1964 4924 2028 4928
rect 1964 4868 1968 4924
rect 1968 4868 2024 4924
rect 2024 4868 2028 4924
rect 1964 4864 2028 4868
rect 2044 4924 2108 4928
rect 2044 4868 2048 4924
rect 2048 4868 2104 4924
rect 2104 4868 2108 4924
rect 2044 4864 2108 4868
rect 2124 4924 2188 4928
rect 2124 4868 2128 4924
rect 2128 4868 2184 4924
rect 2184 4868 2188 4924
rect 2124 4864 2188 4868
rect 2204 4924 2268 4928
rect 2204 4868 2208 4924
rect 2208 4868 2264 4924
rect 2264 4868 2268 4924
rect 2204 4864 2268 4868
rect 3988 4924 4052 4928
rect 3988 4868 3992 4924
rect 3992 4868 4048 4924
rect 4048 4868 4052 4924
rect 3988 4864 4052 4868
rect 4068 4924 4132 4928
rect 4068 4868 4072 4924
rect 4072 4868 4128 4924
rect 4128 4868 4132 4924
rect 4068 4864 4132 4868
rect 4148 4924 4212 4928
rect 4148 4868 4152 4924
rect 4152 4868 4208 4924
rect 4208 4868 4212 4924
rect 4148 4864 4212 4868
rect 4228 4924 4292 4928
rect 4228 4868 4232 4924
rect 4232 4868 4288 4924
rect 4288 4868 4292 4924
rect 4228 4864 4292 4868
rect 6012 4924 6076 4928
rect 6012 4868 6016 4924
rect 6016 4868 6072 4924
rect 6072 4868 6076 4924
rect 6012 4864 6076 4868
rect 6092 4924 6156 4928
rect 6092 4868 6096 4924
rect 6096 4868 6152 4924
rect 6152 4868 6156 4924
rect 6092 4864 6156 4868
rect 6172 4924 6236 4928
rect 6172 4868 6176 4924
rect 6176 4868 6232 4924
rect 6232 4868 6236 4924
rect 6172 4864 6236 4868
rect 6252 4924 6316 4928
rect 6252 4868 6256 4924
rect 6256 4868 6312 4924
rect 6312 4868 6316 4924
rect 6252 4864 6316 4868
rect 8036 4924 8100 4928
rect 8036 4868 8040 4924
rect 8040 4868 8096 4924
rect 8096 4868 8100 4924
rect 8036 4864 8100 4868
rect 8116 4924 8180 4928
rect 8116 4868 8120 4924
rect 8120 4868 8176 4924
rect 8176 4868 8180 4924
rect 8116 4864 8180 4868
rect 8196 4924 8260 4928
rect 8196 4868 8200 4924
rect 8200 4868 8256 4924
rect 8256 4868 8260 4924
rect 8196 4864 8260 4868
rect 8276 4924 8340 4928
rect 8276 4868 8280 4924
rect 8280 4868 8336 4924
rect 8336 4868 8340 4924
rect 8276 4864 8340 4868
rect 2624 4380 2688 4384
rect 2624 4324 2628 4380
rect 2628 4324 2684 4380
rect 2684 4324 2688 4380
rect 2624 4320 2688 4324
rect 2704 4380 2768 4384
rect 2704 4324 2708 4380
rect 2708 4324 2764 4380
rect 2764 4324 2768 4380
rect 2704 4320 2768 4324
rect 2784 4380 2848 4384
rect 2784 4324 2788 4380
rect 2788 4324 2844 4380
rect 2844 4324 2848 4380
rect 2784 4320 2848 4324
rect 2864 4380 2928 4384
rect 2864 4324 2868 4380
rect 2868 4324 2924 4380
rect 2924 4324 2928 4380
rect 2864 4320 2928 4324
rect 4648 4380 4712 4384
rect 4648 4324 4652 4380
rect 4652 4324 4708 4380
rect 4708 4324 4712 4380
rect 4648 4320 4712 4324
rect 4728 4380 4792 4384
rect 4728 4324 4732 4380
rect 4732 4324 4788 4380
rect 4788 4324 4792 4380
rect 4728 4320 4792 4324
rect 4808 4380 4872 4384
rect 4808 4324 4812 4380
rect 4812 4324 4868 4380
rect 4868 4324 4872 4380
rect 4808 4320 4872 4324
rect 4888 4380 4952 4384
rect 4888 4324 4892 4380
rect 4892 4324 4948 4380
rect 4948 4324 4952 4380
rect 4888 4320 4952 4324
rect 6672 4380 6736 4384
rect 6672 4324 6676 4380
rect 6676 4324 6732 4380
rect 6732 4324 6736 4380
rect 6672 4320 6736 4324
rect 6752 4380 6816 4384
rect 6752 4324 6756 4380
rect 6756 4324 6812 4380
rect 6812 4324 6816 4380
rect 6752 4320 6816 4324
rect 6832 4380 6896 4384
rect 6832 4324 6836 4380
rect 6836 4324 6892 4380
rect 6892 4324 6896 4380
rect 6832 4320 6896 4324
rect 6912 4380 6976 4384
rect 6912 4324 6916 4380
rect 6916 4324 6972 4380
rect 6972 4324 6976 4380
rect 6912 4320 6976 4324
rect 8696 4380 8760 4384
rect 8696 4324 8700 4380
rect 8700 4324 8756 4380
rect 8756 4324 8760 4380
rect 8696 4320 8760 4324
rect 8776 4380 8840 4384
rect 8776 4324 8780 4380
rect 8780 4324 8836 4380
rect 8836 4324 8840 4380
rect 8776 4320 8840 4324
rect 8856 4380 8920 4384
rect 8856 4324 8860 4380
rect 8860 4324 8916 4380
rect 8916 4324 8920 4380
rect 8856 4320 8920 4324
rect 8936 4380 9000 4384
rect 8936 4324 8940 4380
rect 8940 4324 8996 4380
rect 8996 4324 9000 4380
rect 8936 4320 9000 4324
rect 1964 3836 2028 3840
rect 1964 3780 1968 3836
rect 1968 3780 2024 3836
rect 2024 3780 2028 3836
rect 1964 3776 2028 3780
rect 2044 3836 2108 3840
rect 2044 3780 2048 3836
rect 2048 3780 2104 3836
rect 2104 3780 2108 3836
rect 2044 3776 2108 3780
rect 2124 3836 2188 3840
rect 2124 3780 2128 3836
rect 2128 3780 2184 3836
rect 2184 3780 2188 3836
rect 2124 3776 2188 3780
rect 2204 3836 2268 3840
rect 2204 3780 2208 3836
rect 2208 3780 2264 3836
rect 2264 3780 2268 3836
rect 2204 3776 2268 3780
rect 3988 3836 4052 3840
rect 3988 3780 3992 3836
rect 3992 3780 4048 3836
rect 4048 3780 4052 3836
rect 3988 3776 4052 3780
rect 4068 3836 4132 3840
rect 4068 3780 4072 3836
rect 4072 3780 4128 3836
rect 4128 3780 4132 3836
rect 4068 3776 4132 3780
rect 4148 3836 4212 3840
rect 4148 3780 4152 3836
rect 4152 3780 4208 3836
rect 4208 3780 4212 3836
rect 4148 3776 4212 3780
rect 4228 3836 4292 3840
rect 4228 3780 4232 3836
rect 4232 3780 4288 3836
rect 4288 3780 4292 3836
rect 4228 3776 4292 3780
rect 6012 3836 6076 3840
rect 6012 3780 6016 3836
rect 6016 3780 6072 3836
rect 6072 3780 6076 3836
rect 6012 3776 6076 3780
rect 6092 3836 6156 3840
rect 6092 3780 6096 3836
rect 6096 3780 6152 3836
rect 6152 3780 6156 3836
rect 6092 3776 6156 3780
rect 6172 3836 6236 3840
rect 6172 3780 6176 3836
rect 6176 3780 6232 3836
rect 6232 3780 6236 3836
rect 6172 3776 6236 3780
rect 6252 3836 6316 3840
rect 6252 3780 6256 3836
rect 6256 3780 6312 3836
rect 6312 3780 6316 3836
rect 6252 3776 6316 3780
rect 8036 3836 8100 3840
rect 8036 3780 8040 3836
rect 8040 3780 8096 3836
rect 8096 3780 8100 3836
rect 8036 3776 8100 3780
rect 8116 3836 8180 3840
rect 8116 3780 8120 3836
rect 8120 3780 8176 3836
rect 8176 3780 8180 3836
rect 8116 3776 8180 3780
rect 8196 3836 8260 3840
rect 8196 3780 8200 3836
rect 8200 3780 8256 3836
rect 8256 3780 8260 3836
rect 8196 3776 8260 3780
rect 8276 3836 8340 3840
rect 8276 3780 8280 3836
rect 8280 3780 8336 3836
rect 8336 3780 8340 3836
rect 8276 3776 8340 3780
rect 2624 3292 2688 3296
rect 2624 3236 2628 3292
rect 2628 3236 2684 3292
rect 2684 3236 2688 3292
rect 2624 3232 2688 3236
rect 2704 3292 2768 3296
rect 2704 3236 2708 3292
rect 2708 3236 2764 3292
rect 2764 3236 2768 3292
rect 2704 3232 2768 3236
rect 2784 3292 2848 3296
rect 2784 3236 2788 3292
rect 2788 3236 2844 3292
rect 2844 3236 2848 3292
rect 2784 3232 2848 3236
rect 2864 3292 2928 3296
rect 2864 3236 2868 3292
rect 2868 3236 2924 3292
rect 2924 3236 2928 3292
rect 2864 3232 2928 3236
rect 4648 3292 4712 3296
rect 4648 3236 4652 3292
rect 4652 3236 4708 3292
rect 4708 3236 4712 3292
rect 4648 3232 4712 3236
rect 4728 3292 4792 3296
rect 4728 3236 4732 3292
rect 4732 3236 4788 3292
rect 4788 3236 4792 3292
rect 4728 3232 4792 3236
rect 4808 3292 4872 3296
rect 4808 3236 4812 3292
rect 4812 3236 4868 3292
rect 4868 3236 4872 3292
rect 4808 3232 4872 3236
rect 4888 3292 4952 3296
rect 4888 3236 4892 3292
rect 4892 3236 4948 3292
rect 4948 3236 4952 3292
rect 4888 3232 4952 3236
rect 6672 3292 6736 3296
rect 6672 3236 6676 3292
rect 6676 3236 6732 3292
rect 6732 3236 6736 3292
rect 6672 3232 6736 3236
rect 6752 3292 6816 3296
rect 6752 3236 6756 3292
rect 6756 3236 6812 3292
rect 6812 3236 6816 3292
rect 6752 3232 6816 3236
rect 6832 3292 6896 3296
rect 6832 3236 6836 3292
rect 6836 3236 6892 3292
rect 6892 3236 6896 3292
rect 6832 3232 6896 3236
rect 6912 3292 6976 3296
rect 6912 3236 6916 3292
rect 6916 3236 6972 3292
rect 6972 3236 6976 3292
rect 6912 3232 6976 3236
rect 8696 3292 8760 3296
rect 8696 3236 8700 3292
rect 8700 3236 8756 3292
rect 8756 3236 8760 3292
rect 8696 3232 8760 3236
rect 8776 3292 8840 3296
rect 8776 3236 8780 3292
rect 8780 3236 8836 3292
rect 8836 3236 8840 3292
rect 8776 3232 8840 3236
rect 8856 3292 8920 3296
rect 8856 3236 8860 3292
rect 8860 3236 8916 3292
rect 8916 3236 8920 3292
rect 8856 3232 8920 3236
rect 8936 3292 9000 3296
rect 8936 3236 8940 3292
rect 8940 3236 8996 3292
rect 8996 3236 9000 3292
rect 8936 3232 9000 3236
rect 1964 2748 2028 2752
rect 1964 2692 1968 2748
rect 1968 2692 2024 2748
rect 2024 2692 2028 2748
rect 1964 2688 2028 2692
rect 2044 2748 2108 2752
rect 2044 2692 2048 2748
rect 2048 2692 2104 2748
rect 2104 2692 2108 2748
rect 2044 2688 2108 2692
rect 2124 2748 2188 2752
rect 2124 2692 2128 2748
rect 2128 2692 2184 2748
rect 2184 2692 2188 2748
rect 2124 2688 2188 2692
rect 2204 2748 2268 2752
rect 2204 2692 2208 2748
rect 2208 2692 2264 2748
rect 2264 2692 2268 2748
rect 2204 2688 2268 2692
rect 3988 2748 4052 2752
rect 3988 2692 3992 2748
rect 3992 2692 4048 2748
rect 4048 2692 4052 2748
rect 3988 2688 4052 2692
rect 4068 2748 4132 2752
rect 4068 2692 4072 2748
rect 4072 2692 4128 2748
rect 4128 2692 4132 2748
rect 4068 2688 4132 2692
rect 4148 2748 4212 2752
rect 4148 2692 4152 2748
rect 4152 2692 4208 2748
rect 4208 2692 4212 2748
rect 4148 2688 4212 2692
rect 4228 2748 4292 2752
rect 4228 2692 4232 2748
rect 4232 2692 4288 2748
rect 4288 2692 4292 2748
rect 4228 2688 4292 2692
rect 6012 2748 6076 2752
rect 6012 2692 6016 2748
rect 6016 2692 6072 2748
rect 6072 2692 6076 2748
rect 6012 2688 6076 2692
rect 6092 2748 6156 2752
rect 6092 2692 6096 2748
rect 6096 2692 6152 2748
rect 6152 2692 6156 2748
rect 6092 2688 6156 2692
rect 6172 2748 6236 2752
rect 6172 2692 6176 2748
rect 6176 2692 6232 2748
rect 6232 2692 6236 2748
rect 6172 2688 6236 2692
rect 6252 2748 6316 2752
rect 6252 2692 6256 2748
rect 6256 2692 6312 2748
rect 6312 2692 6316 2748
rect 6252 2688 6316 2692
rect 8036 2748 8100 2752
rect 8036 2692 8040 2748
rect 8040 2692 8096 2748
rect 8096 2692 8100 2748
rect 8036 2688 8100 2692
rect 8116 2748 8180 2752
rect 8116 2692 8120 2748
rect 8120 2692 8176 2748
rect 8176 2692 8180 2748
rect 8116 2688 8180 2692
rect 8196 2748 8260 2752
rect 8196 2692 8200 2748
rect 8200 2692 8256 2748
rect 8256 2692 8260 2748
rect 8196 2688 8260 2692
rect 8276 2748 8340 2752
rect 8276 2692 8280 2748
rect 8280 2692 8336 2748
rect 8336 2692 8340 2748
rect 8276 2688 8340 2692
rect 2624 2204 2688 2208
rect 2624 2148 2628 2204
rect 2628 2148 2684 2204
rect 2684 2148 2688 2204
rect 2624 2144 2688 2148
rect 2704 2204 2768 2208
rect 2704 2148 2708 2204
rect 2708 2148 2764 2204
rect 2764 2148 2768 2204
rect 2704 2144 2768 2148
rect 2784 2204 2848 2208
rect 2784 2148 2788 2204
rect 2788 2148 2844 2204
rect 2844 2148 2848 2204
rect 2784 2144 2848 2148
rect 2864 2204 2928 2208
rect 2864 2148 2868 2204
rect 2868 2148 2924 2204
rect 2924 2148 2928 2204
rect 2864 2144 2928 2148
rect 4648 2204 4712 2208
rect 4648 2148 4652 2204
rect 4652 2148 4708 2204
rect 4708 2148 4712 2204
rect 4648 2144 4712 2148
rect 4728 2204 4792 2208
rect 4728 2148 4732 2204
rect 4732 2148 4788 2204
rect 4788 2148 4792 2204
rect 4728 2144 4792 2148
rect 4808 2204 4872 2208
rect 4808 2148 4812 2204
rect 4812 2148 4868 2204
rect 4868 2148 4872 2204
rect 4808 2144 4872 2148
rect 4888 2204 4952 2208
rect 4888 2148 4892 2204
rect 4892 2148 4948 2204
rect 4948 2148 4952 2204
rect 4888 2144 4952 2148
rect 6672 2204 6736 2208
rect 6672 2148 6676 2204
rect 6676 2148 6732 2204
rect 6732 2148 6736 2204
rect 6672 2144 6736 2148
rect 6752 2204 6816 2208
rect 6752 2148 6756 2204
rect 6756 2148 6812 2204
rect 6812 2148 6816 2204
rect 6752 2144 6816 2148
rect 6832 2204 6896 2208
rect 6832 2148 6836 2204
rect 6836 2148 6892 2204
rect 6892 2148 6896 2204
rect 6832 2144 6896 2148
rect 6912 2204 6976 2208
rect 6912 2148 6916 2204
rect 6916 2148 6972 2204
rect 6972 2148 6976 2204
rect 6912 2144 6976 2148
rect 8696 2204 8760 2208
rect 8696 2148 8700 2204
rect 8700 2148 8756 2204
rect 8756 2148 8760 2204
rect 8696 2144 8760 2148
rect 8776 2204 8840 2208
rect 8776 2148 8780 2204
rect 8780 2148 8836 2204
rect 8836 2148 8840 2204
rect 8776 2144 8840 2148
rect 8856 2204 8920 2208
rect 8856 2148 8860 2204
rect 8860 2148 8916 2204
rect 8916 2148 8920 2204
rect 8856 2144 8920 2148
rect 8936 2204 9000 2208
rect 8936 2148 8940 2204
rect 8940 2148 8996 2204
rect 8996 2148 9000 2204
rect 8936 2144 9000 2148
<< metal4 >>
rect 1956 9280 2276 9840
rect 1956 9216 1964 9280
rect 2028 9216 2044 9280
rect 2108 9216 2124 9280
rect 2188 9216 2204 9280
rect 2268 9216 2276 9280
rect 1956 8958 2276 9216
rect 1956 8722 1998 8958
rect 2234 8722 2276 8958
rect 1956 8192 2276 8722
rect 1956 8128 1964 8192
rect 2028 8128 2044 8192
rect 2108 8128 2124 8192
rect 2188 8128 2204 8192
rect 2268 8128 2276 8192
rect 1956 7104 2276 8128
rect 1956 7040 1964 7104
rect 2028 7054 2044 7104
rect 2108 7054 2124 7104
rect 2188 7054 2204 7104
rect 2268 7040 2276 7104
rect 1956 6818 1998 7040
rect 2234 6818 2276 7040
rect 1956 6016 2276 6818
rect 1956 5952 1964 6016
rect 2028 5952 2044 6016
rect 2108 5952 2124 6016
rect 2188 5952 2204 6016
rect 2268 5952 2276 6016
rect 1956 5150 2276 5952
rect 1956 4928 1998 5150
rect 2234 4928 2276 5150
rect 1956 4864 1964 4928
rect 2028 4864 2044 4914
rect 2108 4864 2124 4914
rect 2188 4864 2204 4914
rect 2268 4864 2276 4928
rect 1956 3840 2276 4864
rect 1956 3776 1964 3840
rect 2028 3776 2044 3840
rect 2108 3776 2124 3840
rect 2188 3776 2204 3840
rect 2268 3776 2276 3840
rect 1956 3246 2276 3776
rect 1956 3010 1998 3246
rect 2234 3010 2276 3246
rect 1956 2752 2276 3010
rect 1956 2688 1964 2752
rect 2028 2688 2044 2752
rect 2108 2688 2124 2752
rect 2188 2688 2204 2752
rect 2268 2688 2276 2752
rect 1956 2128 2276 2688
rect 2616 9824 2936 9840
rect 2616 9760 2624 9824
rect 2688 9760 2704 9824
rect 2768 9760 2784 9824
rect 2848 9760 2864 9824
rect 2928 9760 2936 9824
rect 2616 9618 2936 9760
rect 2616 9382 2658 9618
rect 2894 9382 2936 9618
rect 2616 8736 2936 9382
rect 2616 8672 2624 8736
rect 2688 8672 2704 8736
rect 2768 8672 2784 8736
rect 2848 8672 2864 8736
rect 2928 8672 2936 8736
rect 2616 7714 2936 8672
rect 2616 7648 2658 7714
rect 2894 7648 2936 7714
rect 2616 7584 2624 7648
rect 2928 7584 2936 7648
rect 2616 7478 2658 7584
rect 2894 7478 2936 7584
rect 2616 6560 2936 7478
rect 2616 6496 2624 6560
rect 2688 6496 2704 6560
rect 2768 6496 2784 6560
rect 2848 6496 2864 6560
rect 2928 6496 2936 6560
rect 2616 5810 2936 6496
rect 2616 5574 2658 5810
rect 2894 5574 2936 5810
rect 2616 5472 2936 5574
rect 2616 5408 2624 5472
rect 2688 5408 2704 5472
rect 2768 5408 2784 5472
rect 2848 5408 2864 5472
rect 2928 5408 2936 5472
rect 2616 4384 2936 5408
rect 2616 4320 2624 4384
rect 2688 4320 2704 4384
rect 2768 4320 2784 4384
rect 2848 4320 2864 4384
rect 2928 4320 2936 4384
rect 2616 3906 2936 4320
rect 2616 3670 2658 3906
rect 2894 3670 2936 3906
rect 2616 3296 2936 3670
rect 2616 3232 2624 3296
rect 2688 3232 2704 3296
rect 2768 3232 2784 3296
rect 2848 3232 2864 3296
rect 2928 3232 2936 3296
rect 2616 2208 2936 3232
rect 2616 2144 2624 2208
rect 2688 2144 2704 2208
rect 2768 2144 2784 2208
rect 2848 2144 2864 2208
rect 2928 2144 2936 2208
rect 2616 2128 2936 2144
rect 3980 9280 4300 9840
rect 3980 9216 3988 9280
rect 4052 9216 4068 9280
rect 4132 9216 4148 9280
rect 4212 9216 4228 9280
rect 4292 9216 4300 9280
rect 3980 8958 4300 9216
rect 3980 8722 4022 8958
rect 4258 8722 4300 8958
rect 3980 8192 4300 8722
rect 3980 8128 3988 8192
rect 4052 8128 4068 8192
rect 4132 8128 4148 8192
rect 4212 8128 4228 8192
rect 4292 8128 4300 8192
rect 3980 7104 4300 8128
rect 3980 7040 3988 7104
rect 4052 7054 4068 7104
rect 4132 7054 4148 7104
rect 4212 7054 4228 7104
rect 4292 7040 4300 7104
rect 3980 6818 4022 7040
rect 4258 6818 4300 7040
rect 3980 6016 4300 6818
rect 3980 5952 3988 6016
rect 4052 5952 4068 6016
rect 4132 5952 4148 6016
rect 4212 5952 4228 6016
rect 4292 5952 4300 6016
rect 3980 5150 4300 5952
rect 3980 4928 4022 5150
rect 4258 4928 4300 5150
rect 3980 4864 3988 4928
rect 4052 4864 4068 4914
rect 4132 4864 4148 4914
rect 4212 4864 4228 4914
rect 4292 4864 4300 4928
rect 3980 3840 4300 4864
rect 3980 3776 3988 3840
rect 4052 3776 4068 3840
rect 4132 3776 4148 3840
rect 4212 3776 4228 3840
rect 4292 3776 4300 3840
rect 3980 3246 4300 3776
rect 3980 3010 4022 3246
rect 4258 3010 4300 3246
rect 3980 2752 4300 3010
rect 3980 2688 3988 2752
rect 4052 2688 4068 2752
rect 4132 2688 4148 2752
rect 4212 2688 4228 2752
rect 4292 2688 4300 2752
rect 3980 2128 4300 2688
rect 4640 9824 4960 9840
rect 4640 9760 4648 9824
rect 4712 9760 4728 9824
rect 4792 9760 4808 9824
rect 4872 9760 4888 9824
rect 4952 9760 4960 9824
rect 4640 9618 4960 9760
rect 4640 9382 4682 9618
rect 4918 9382 4960 9618
rect 4640 8736 4960 9382
rect 4640 8672 4648 8736
rect 4712 8672 4728 8736
rect 4792 8672 4808 8736
rect 4872 8672 4888 8736
rect 4952 8672 4960 8736
rect 4640 7714 4960 8672
rect 4640 7648 4682 7714
rect 4918 7648 4960 7714
rect 4640 7584 4648 7648
rect 4952 7584 4960 7648
rect 4640 7478 4682 7584
rect 4918 7478 4960 7584
rect 4640 6560 4960 7478
rect 4640 6496 4648 6560
rect 4712 6496 4728 6560
rect 4792 6496 4808 6560
rect 4872 6496 4888 6560
rect 4952 6496 4960 6560
rect 4640 5810 4960 6496
rect 4640 5574 4682 5810
rect 4918 5574 4960 5810
rect 4640 5472 4960 5574
rect 4640 5408 4648 5472
rect 4712 5408 4728 5472
rect 4792 5408 4808 5472
rect 4872 5408 4888 5472
rect 4952 5408 4960 5472
rect 4640 4384 4960 5408
rect 4640 4320 4648 4384
rect 4712 4320 4728 4384
rect 4792 4320 4808 4384
rect 4872 4320 4888 4384
rect 4952 4320 4960 4384
rect 4640 3906 4960 4320
rect 4640 3670 4682 3906
rect 4918 3670 4960 3906
rect 4640 3296 4960 3670
rect 4640 3232 4648 3296
rect 4712 3232 4728 3296
rect 4792 3232 4808 3296
rect 4872 3232 4888 3296
rect 4952 3232 4960 3296
rect 4640 2208 4960 3232
rect 4640 2144 4648 2208
rect 4712 2144 4728 2208
rect 4792 2144 4808 2208
rect 4872 2144 4888 2208
rect 4952 2144 4960 2208
rect 4640 2128 4960 2144
rect 6004 9280 6324 9840
rect 6004 9216 6012 9280
rect 6076 9216 6092 9280
rect 6156 9216 6172 9280
rect 6236 9216 6252 9280
rect 6316 9216 6324 9280
rect 6004 8958 6324 9216
rect 6004 8722 6046 8958
rect 6282 8722 6324 8958
rect 6004 8192 6324 8722
rect 6004 8128 6012 8192
rect 6076 8128 6092 8192
rect 6156 8128 6172 8192
rect 6236 8128 6252 8192
rect 6316 8128 6324 8192
rect 6004 7104 6324 8128
rect 6004 7040 6012 7104
rect 6076 7054 6092 7104
rect 6156 7054 6172 7104
rect 6236 7054 6252 7104
rect 6316 7040 6324 7104
rect 6004 6818 6046 7040
rect 6282 6818 6324 7040
rect 6004 6016 6324 6818
rect 6004 5952 6012 6016
rect 6076 5952 6092 6016
rect 6156 5952 6172 6016
rect 6236 5952 6252 6016
rect 6316 5952 6324 6016
rect 6004 5150 6324 5952
rect 6004 4928 6046 5150
rect 6282 4928 6324 5150
rect 6004 4864 6012 4928
rect 6076 4864 6092 4914
rect 6156 4864 6172 4914
rect 6236 4864 6252 4914
rect 6316 4864 6324 4928
rect 6004 3840 6324 4864
rect 6004 3776 6012 3840
rect 6076 3776 6092 3840
rect 6156 3776 6172 3840
rect 6236 3776 6252 3840
rect 6316 3776 6324 3840
rect 6004 3246 6324 3776
rect 6004 3010 6046 3246
rect 6282 3010 6324 3246
rect 6004 2752 6324 3010
rect 6004 2688 6012 2752
rect 6076 2688 6092 2752
rect 6156 2688 6172 2752
rect 6236 2688 6252 2752
rect 6316 2688 6324 2752
rect 6004 2128 6324 2688
rect 6664 9824 6984 9840
rect 6664 9760 6672 9824
rect 6736 9760 6752 9824
rect 6816 9760 6832 9824
rect 6896 9760 6912 9824
rect 6976 9760 6984 9824
rect 6664 9618 6984 9760
rect 6664 9382 6706 9618
rect 6942 9382 6984 9618
rect 6664 8736 6984 9382
rect 6664 8672 6672 8736
rect 6736 8672 6752 8736
rect 6816 8672 6832 8736
rect 6896 8672 6912 8736
rect 6976 8672 6984 8736
rect 6664 7714 6984 8672
rect 6664 7648 6706 7714
rect 6942 7648 6984 7714
rect 6664 7584 6672 7648
rect 6976 7584 6984 7648
rect 6664 7478 6706 7584
rect 6942 7478 6984 7584
rect 6664 6560 6984 7478
rect 6664 6496 6672 6560
rect 6736 6496 6752 6560
rect 6816 6496 6832 6560
rect 6896 6496 6912 6560
rect 6976 6496 6984 6560
rect 6664 5810 6984 6496
rect 6664 5574 6706 5810
rect 6942 5574 6984 5810
rect 6664 5472 6984 5574
rect 6664 5408 6672 5472
rect 6736 5408 6752 5472
rect 6816 5408 6832 5472
rect 6896 5408 6912 5472
rect 6976 5408 6984 5472
rect 6664 4384 6984 5408
rect 6664 4320 6672 4384
rect 6736 4320 6752 4384
rect 6816 4320 6832 4384
rect 6896 4320 6912 4384
rect 6976 4320 6984 4384
rect 6664 3906 6984 4320
rect 6664 3670 6706 3906
rect 6942 3670 6984 3906
rect 6664 3296 6984 3670
rect 6664 3232 6672 3296
rect 6736 3232 6752 3296
rect 6816 3232 6832 3296
rect 6896 3232 6912 3296
rect 6976 3232 6984 3296
rect 6664 2208 6984 3232
rect 6664 2144 6672 2208
rect 6736 2144 6752 2208
rect 6816 2144 6832 2208
rect 6896 2144 6912 2208
rect 6976 2144 6984 2208
rect 6664 2128 6984 2144
rect 8028 9280 8348 9840
rect 8028 9216 8036 9280
rect 8100 9216 8116 9280
rect 8180 9216 8196 9280
rect 8260 9216 8276 9280
rect 8340 9216 8348 9280
rect 8028 8958 8348 9216
rect 8028 8722 8070 8958
rect 8306 8722 8348 8958
rect 8028 8192 8348 8722
rect 8028 8128 8036 8192
rect 8100 8128 8116 8192
rect 8180 8128 8196 8192
rect 8260 8128 8276 8192
rect 8340 8128 8348 8192
rect 8028 7104 8348 8128
rect 8028 7040 8036 7104
rect 8100 7054 8116 7104
rect 8180 7054 8196 7104
rect 8260 7054 8276 7104
rect 8340 7040 8348 7104
rect 8028 6818 8070 7040
rect 8306 6818 8348 7040
rect 8028 6016 8348 6818
rect 8028 5952 8036 6016
rect 8100 5952 8116 6016
rect 8180 5952 8196 6016
rect 8260 5952 8276 6016
rect 8340 5952 8348 6016
rect 8028 5150 8348 5952
rect 8028 4928 8070 5150
rect 8306 4928 8348 5150
rect 8028 4864 8036 4928
rect 8100 4864 8116 4914
rect 8180 4864 8196 4914
rect 8260 4864 8276 4914
rect 8340 4864 8348 4928
rect 8028 3840 8348 4864
rect 8028 3776 8036 3840
rect 8100 3776 8116 3840
rect 8180 3776 8196 3840
rect 8260 3776 8276 3840
rect 8340 3776 8348 3840
rect 8028 3246 8348 3776
rect 8028 3010 8070 3246
rect 8306 3010 8348 3246
rect 8028 2752 8348 3010
rect 8028 2688 8036 2752
rect 8100 2688 8116 2752
rect 8180 2688 8196 2752
rect 8260 2688 8276 2752
rect 8340 2688 8348 2752
rect 8028 2128 8348 2688
rect 8688 9824 9008 9840
rect 8688 9760 8696 9824
rect 8760 9760 8776 9824
rect 8840 9760 8856 9824
rect 8920 9760 8936 9824
rect 9000 9760 9008 9824
rect 8688 9618 9008 9760
rect 8688 9382 8730 9618
rect 8966 9382 9008 9618
rect 8688 8736 9008 9382
rect 8688 8672 8696 8736
rect 8760 8672 8776 8736
rect 8840 8672 8856 8736
rect 8920 8672 8936 8736
rect 9000 8672 9008 8736
rect 8688 7714 9008 8672
rect 8688 7648 8730 7714
rect 8966 7648 9008 7714
rect 8688 7584 8696 7648
rect 9000 7584 9008 7648
rect 8688 7478 8730 7584
rect 8966 7478 9008 7584
rect 8688 6560 9008 7478
rect 8688 6496 8696 6560
rect 8760 6496 8776 6560
rect 8840 6496 8856 6560
rect 8920 6496 8936 6560
rect 9000 6496 9008 6560
rect 8688 5810 9008 6496
rect 8688 5574 8730 5810
rect 8966 5574 9008 5810
rect 8688 5472 9008 5574
rect 8688 5408 8696 5472
rect 8760 5408 8776 5472
rect 8840 5408 8856 5472
rect 8920 5408 8936 5472
rect 9000 5408 9008 5472
rect 8688 4384 9008 5408
rect 8688 4320 8696 4384
rect 8760 4320 8776 4384
rect 8840 4320 8856 4384
rect 8920 4320 8936 4384
rect 9000 4320 9008 4384
rect 8688 3906 9008 4320
rect 8688 3670 8730 3906
rect 8966 3670 9008 3906
rect 8688 3296 9008 3670
rect 8688 3232 8696 3296
rect 8760 3232 8776 3296
rect 8840 3232 8856 3296
rect 8920 3232 8936 3296
rect 9000 3232 9008 3296
rect 8688 2208 9008 3232
rect 8688 2144 8696 2208
rect 8760 2144 8776 2208
rect 8840 2144 8856 2208
rect 8920 2144 8936 2208
rect 9000 2144 9008 2208
rect 8688 2128 9008 2144
<< via4 >>
rect 1998 8722 2234 8958
rect 1998 7040 2028 7054
rect 2028 7040 2044 7054
rect 2044 7040 2108 7054
rect 2108 7040 2124 7054
rect 2124 7040 2188 7054
rect 2188 7040 2204 7054
rect 2204 7040 2234 7054
rect 1998 6818 2234 7040
rect 1998 4928 2234 5150
rect 1998 4914 2028 4928
rect 2028 4914 2044 4928
rect 2044 4914 2108 4928
rect 2108 4914 2124 4928
rect 2124 4914 2188 4928
rect 2188 4914 2204 4928
rect 2204 4914 2234 4928
rect 1998 3010 2234 3246
rect 2658 9382 2894 9618
rect 2658 7648 2894 7714
rect 2658 7584 2688 7648
rect 2688 7584 2704 7648
rect 2704 7584 2768 7648
rect 2768 7584 2784 7648
rect 2784 7584 2848 7648
rect 2848 7584 2864 7648
rect 2864 7584 2894 7648
rect 2658 7478 2894 7584
rect 2658 5574 2894 5810
rect 2658 3670 2894 3906
rect 4022 8722 4258 8958
rect 4022 7040 4052 7054
rect 4052 7040 4068 7054
rect 4068 7040 4132 7054
rect 4132 7040 4148 7054
rect 4148 7040 4212 7054
rect 4212 7040 4228 7054
rect 4228 7040 4258 7054
rect 4022 6818 4258 7040
rect 4022 4928 4258 5150
rect 4022 4914 4052 4928
rect 4052 4914 4068 4928
rect 4068 4914 4132 4928
rect 4132 4914 4148 4928
rect 4148 4914 4212 4928
rect 4212 4914 4228 4928
rect 4228 4914 4258 4928
rect 4022 3010 4258 3246
rect 4682 9382 4918 9618
rect 4682 7648 4918 7714
rect 4682 7584 4712 7648
rect 4712 7584 4728 7648
rect 4728 7584 4792 7648
rect 4792 7584 4808 7648
rect 4808 7584 4872 7648
rect 4872 7584 4888 7648
rect 4888 7584 4918 7648
rect 4682 7478 4918 7584
rect 4682 5574 4918 5810
rect 4682 3670 4918 3906
rect 6046 8722 6282 8958
rect 6046 7040 6076 7054
rect 6076 7040 6092 7054
rect 6092 7040 6156 7054
rect 6156 7040 6172 7054
rect 6172 7040 6236 7054
rect 6236 7040 6252 7054
rect 6252 7040 6282 7054
rect 6046 6818 6282 7040
rect 6046 4928 6282 5150
rect 6046 4914 6076 4928
rect 6076 4914 6092 4928
rect 6092 4914 6156 4928
rect 6156 4914 6172 4928
rect 6172 4914 6236 4928
rect 6236 4914 6252 4928
rect 6252 4914 6282 4928
rect 6046 3010 6282 3246
rect 6706 9382 6942 9618
rect 6706 7648 6942 7714
rect 6706 7584 6736 7648
rect 6736 7584 6752 7648
rect 6752 7584 6816 7648
rect 6816 7584 6832 7648
rect 6832 7584 6896 7648
rect 6896 7584 6912 7648
rect 6912 7584 6942 7648
rect 6706 7478 6942 7584
rect 6706 5574 6942 5810
rect 6706 3670 6942 3906
rect 8070 8722 8306 8958
rect 8070 7040 8100 7054
rect 8100 7040 8116 7054
rect 8116 7040 8180 7054
rect 8180 7040 8196 7054
rect 8196 7040 8260 7054
rect 8260 7040 8276 7054
rect 8276 7040 8306 7054
rect 8070 6818 8306 7040
rect 8070 4928 8306 5150
rect 8070 4914 8100 4928
rect 8100 4914 8116 4928
rect 8116 4914 8180 4928
rect 8180 4914 8196 4928
rect 8196 4914 8260 4928
rect 8260 4914 8276 4928
rect 8276 4914 8306 4928
rect 8070 3010 8306 3246
rect 8730 9382 8966 9618
rect 8730 7648 8966 7714
rect 8730 7584 8760 7648
rect 8760 7584 8776 7648
rect 8776 7584 8840 7648
rect 8840 7584 8856 7648
rect 8856 7584 8920 7648
rect 8920 7584 8936 7648
rect 8936 7584 8966 7648
rect 8730 7478 8966 7584
rect 8730 5574 8966 5810
rect 8730 3670 8966 3906
<< metal5 >>
rect 1056 9618 9248 9660
rect 1056 9382 2658 9618
rect 2894 9382 4682 9618
rect 4918 9382 6706 9618
rect 6942 9382 8730 9618
rect 8966 9382 9248 9618
rect 1056 9340 9248 9382
rect 1056 8958 9248 9000
rect 1056 8722 1998 8958
rect 2234 8722 4022 8958
rect 4258 8722 6046 8958
rect 6282 8722 8070 8958
rect 8306 8722 9248 8958
rect 1056 8680 9248 8722
rect 1056 7714 9248 7756
rect 1056 7478 2658 7714
rect 2894 7478 4682 7714
rect 4918 7478 6706 7714
rect 6942 7478 8730 7714
rect 8966 7478 9248 7714
rect 1056 7436 9248 7478
rect 1056 7054 9248 7096
rect 1056 6818 1998 7054
rect 2234 6818 4022 7054
rect 4258 6818 6046 7054
rect 6282 6818 8070 7054
rect 8306 6818 9248 7054
rect 1056 6776 9248 6818
rect 1056 5810 9248 5852
rect 1056 5574 2658 5810
rect 2894 5574 4682 5810
rect 4918 5574 6706 5810
rect 6942 5574 8730 5810
rect 8966 5574 9248 5810
rect 1056 5532 9248 5574
rect 1056 5150 9248 5192
rect 1056 4914 1998 5150
rect 2234 4914 4022 5150
rect 4258 4914 6046 5150
rect 6282 4914 8070 5150
rect 8306 4914 9248 5150
rect 1056 4872 9248 4914
rect 1056 3906 9248 3948
rect 1056 3670 2658 3906
rect 2894 3670 4682 3906
rect 4918 3670 6706 3906
rect 6942 3670 8730 3906
rect 8966 3670 9248 3906
rect 1056 3628 9248 3670
rect 1056 3246 9248 3288
rect 1056 3010 1998 3246
rect 2234 3010 4022 3246
rect 4258 3010 6046 3246
rect 6282 3010 8070 3246
rect 8306 3010 9248 3246
rect 1056 2968 9248 3010
use sky130_fd_sc_hd__inv_2  _043_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _044_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 7820 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _045_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 8096 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _046_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 8280 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _047_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 7912 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _048_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 7820 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _049_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 8188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _050_
timestamp 1704988097
transform 1 0 7268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _051_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 7544 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _052_
timestamp 1704988097
transform 1 0 7636 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _053_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 7360 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _054_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 8188 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _055_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 7544 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _056_
timestamp 1704988097
transform 1 0 8648 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _057_
timestamp 1704988097
transform 1 0 7544 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _058_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 8464 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _059_
timestamp 1704988097
transform 1 0 7452 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _060_
timestamp 1704988097
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 3956 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _062_
timestamp 1704988097
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 5244 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _064_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 3864 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _065_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 4416 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 4508 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1704988097
transform -1 0 2208 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _068_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 4784 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _069_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 4048 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _070_
timestamp 1704988097
transform -1 0 5152 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _071_
timestamp 1704988097
transform -1 0 5428 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _072_
timestamp 1704988097
transform -1 0 2668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 2024 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _074_
timestamp 1704988097
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o31a_1  _075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 2668 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _076_
timestamp 1704988097
transform 1 0 2852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _077_
timestamp 1704988097
transform 1 0 4140 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _078_
timestamp 1704988097
transform -1 0 6072 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _079_
timestamp 1704988097
transform -1 0 4140 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1704988097
transform 1 0 5704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or4_2  _081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 5888 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _082_
timestamp 1704988097
transform -1 0 3680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _083_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 4048 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _084_
timestamp 1704988097
transform 1 0 2852 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _085_
timestamp 1704988097
transform -1 0 4232 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _086_
timestamp 1704988097
transform -1 0 2852 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _087_
timestamp 1704988097
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _088_
timestamp 1704988097
transform 1 0 3312 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor3_1  _089_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 2944 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _090_
timestamp 1704988097
transform 1 0 1932 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _091_
timestamp 1704988097
transform -1 0 2208 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o41a_1  _092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 2668 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _093_
timestamp 1704988097
transform 1 0 2208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_1  _094_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 4048 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _095_
timestamp 1704988097
transform 1 0 4692 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _096_
timestamp 1704988097
transform 1 0 2208 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _097_
timestamp 1704988097
transform 1 0 4416 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _098_
timestamp 1704988097
transform 1 0 1380 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _099_
timestamp 1704988097
transform 1 0 1932 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _100_
timestamp 1704988097
transform 1 0 4508 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _101_
timestamp 1704988097
transform 1 0 3772 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _102_
timestamp 1704988097
transform 1 0 1380 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _103_
timestamp 1704988097
transform 1 0 1380 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _104_
timestamp 1704988097
transform -1 0 2944 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _105_
timestamp 1704988097
transform 1 0 5888 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _106_
timestamp 1704988097
transform 1 0 6348 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _107_
timestamp 1704988097
transform 1 0 5612 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _108_
timestamp 1704988097
transform 1 0 6348 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _109_
timestamp 1704988097
transform 1 0 5520 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _110_
timestamp 1704988097
transform 1 0 6348 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _111_
timestamp 1704988097
transform 1 0 6348 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _112_
timestamp 1704988097
transform 1 0 5980 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 3772 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1704988097
transform -1 0 4692 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1704988097
transform 1 0 3128 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 1380 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_37
timestamp 1704988097
transform 1 0 4508 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 4968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1704988097
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_69
timestamp 1704988097
transform 1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_77
timestamp 1704988097
transform 1 0 8188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1704988097
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_83
timestamp 1704988097
transform 1 0 8740 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_10
timestamp 1704988097
transform 1 0 2024 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_22
timestamp 1704988097
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_29
timestamp 1704988097
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 4876 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_68
timestamp 1704988097
transform 1 0 7360 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_72
timestamp 1704988097
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_76
timestamp 1704988097
transform 1 0 8096 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 1380 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_11
timestamp 1704988097
transform 1 0 2116 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_19
timestamp 1704988097
transform 1 0 2852 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_31
timestamp 1704988097
transform 1 0 3956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_39
timestamp 1704988097
transform 1 0 4692 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_45
timestamp 1704988097
transform 1 0 5244 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_53
timestamp 1704988097
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1704988097
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_77
timestamp 1704988097
transform 1 0 8188 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_25
timestamp 1704988097
transform 1 0 3404 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_47
timestamp 1704988097
transform 1 0 5428 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_65
timestamp 1704988097
transform 1 0 7084 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_78
timestamp 1704988097
transform 1 0 8280 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_3
timestamp 1704988097
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_29
timestamp 1704988097
transform 1 0 3772 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_34
timestamp 1704988097
transform 1 0 4232 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_52
timestamp 1704988097
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_80
timestamp 1704988097
transform 1 0 8464 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_20
timestamp 1704988097
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_57
timestamp 1704988097
transform 1 0 6348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_69
timestamp 1704988097
transform 1 0 7452 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_74
timestamp 1704988097
transform 1 0 7912 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_3
timestamp 1704988097
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_15
timestamp 1704988097
transform 1 0 2484 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_26
timestamp 1704988097
transform 1 0 3496 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_48
timestamp 1704988097
transform 1 0 5520 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_52
timestamp 1704988097
transform 1 0 5888 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1704988097
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_65
timestamp 1704988097
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_75
timestamp 1704988097
transform 1 0 8004 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1704988097
transform 1 0 1380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_20
timestamp 1704988097
transform 1 0 2944 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_24
timestamp 1704988097
transform 1 0 3312 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_39
timestamp 1704988097
transform 1 0 4692 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_47
timestamp 1704988097
transform 1 0 5428 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_64
timestamp 1704988097
transform 1 0 6992 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_77
timestamp 1704988097
transform 1 0 8188 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_3
timestamp 1704988097
transform 1 0 1380 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_11
timestamp 1704988097
transform 1 0 2116 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_24
timestamp 1704988097
transform 1 0 3312 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_54
timestamp 1704988097
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_80
timestamp 1704988097
transform 1 0 8464 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_84
timestamp 1704988097
transform 1 0 8832 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_7
timestamp 1704988097
transform 1 0 1748 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_52
timestamp 1704988097
transform 1 0 5888 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_64
timestamp 1704988097
transform 1 0 6992 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_76
timestamp 1704988097
transform 1 0 8096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1704988097
transform 1 0 5980 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_73
timestamp 1704988097
transform 1 0 7820 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_3
timestamp 1704988097
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_25
timestamp 1704988097
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_76
timestamp 1704988097
transform 1 0 8096 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1704988097
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1704988097
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_27
timestamp 1704988097
transform 1 0 3588 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_29
timestamp 1704988097
transform 1 0 3772 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_41
timestamp 1704988097
transform 1 0 4876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_53
timestamp 1704988097
transform 1 0 5980 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_61
timestamp 1704988097
transform 1 0 6716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_73
timestamp 1704988097
transform 1 0 7820 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_81
timestamp 1704988097
transform 1 0 8556 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 3312 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  hold2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 6256 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704988097
transform -1 0 6348 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704988097
transform -1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704988097
transform 1 0 1748 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704988097
transform -1 0 5888 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704988097
transform -1 0 5704 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704988097
transform -1 0 4508 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1704988097
transform -1 0 3312 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform -1 0 6716 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1704988097
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 1704988097
transform 1 0 8464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output4 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output5
timestamp 1704988097
transform 1 0 8464 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output6
timestamp 1704988097
transform 1 0 8556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output7
timestamp 1704988097
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output8
timestamp 1704988097
transform -1 0 8832 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output9
timestamp 1704988097
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1704988097
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 1704988097
transform -1 0 1932 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_14
timestamp 1704988097
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704988097
transform -1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_15
timestamp 1704988097
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704988097
transform -1 0 9200 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_16
timestamp 1704988097
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704988097
transform -1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_17
timestamp 1704988097
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704988097
transform -1 0 9200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_18
timestamp 1704988097
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704988097
transform -1 0 9200 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_19
timestamp 1704988097
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704988097
transform -1 0 9200 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_20
timestamp 1704988097
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704988097
transform -1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_21
timestamp 1704988097
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704988097
transform -1 0 9200 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_22
timestamp 1704988097
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704988097
transform -1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_23
timestamp 1704988097
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704988097
transform -1 0 9200 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_24
timestamp 1704988097
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704988097
transform -1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_25
timestamp 1704988097
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704988097
transform -1 0 9200 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_26
timestamp 1704988097
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704988097
transform -1 0 9200 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_27
timestamp 1704988097
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704988097
transform -1 0 9200 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_28 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704988097
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_29
timestamp 1704988097
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_30
timestamp 1704988097
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_31
timestamp 1704988097
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_32
timestamp 1704988097
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_33
timestamp 1704988097
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_34
timestamp 1704988097
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_35
timestamp 1704988097
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_36
timestamp 1704988097
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_37
timestamp 1704988097
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_38
timestamp 1704988097
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_39
timestamp 1704988097
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_40
timestamp 1704988097
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_41
timestamp 1704988097
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_42
timestamp 1704988097
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_43
timestamp 1704988097
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_44
timestamp 1704988097
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_45
timestamp 1704988097
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_46
timestamp 1704988097
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_47
timestamp 1704988097
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_48
timestamp 1704988097
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_49
timestamp 1704988097
transform 1 0 3680 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_50
timestamp 1704988097
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_51
timestamp 1704988097
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
<< labels >>
flabel metal4 s 2616 2128 2936 9840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4640 2128 4960 9840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 6664 2128 6984 9840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 8688 2128 9008 9840 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 3628 9248 3948 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 5532 9248 5852 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 7436 9248 7756 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 9340 9248 9660 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1956 2128 2276 9840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 3980 2128 4300 9840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 6004 2128 6324 9840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 8028 2128 8348 9840 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 2968 9248 3288 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4872 9248 5192 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 6776 9248 7096 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 8680 9248 9000 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 9517 3408 10317 3528 0 FreeSans 480 0 0 0 data_out[0]
port 3 nsew signal tristate
flabel metal3 s 9517 2728 10317 2848 0 FreeSans 480 0 0 0 data_out[1]
port 4 nsew signal tristate
flabel metal3 s 9517 4088 10317 4208 0 FreeSans 480 0 0 0 data_out[2]
port 5 nsew signal tristate
flabel metal3 s 9517 4768 10317 4888 0 FreeSans 480 0 0 0 data_out[3]
port 6 nsew signal tristate
flabel metal3 s 9517 6128 10317 6248 0 FreeSans 480 0 0 0 data_out[4]
port 7 nsew signal tristate
flabel metal3 s 9517 6808 10317 6928 0 FreeSans 480 0 0 0 data_out[5]
port 8 nsew signal tristate
flabel metal3 s 9517 7488 10317 7608 0 FreeSans 480 0 0 0 data_out[6]
port 9 nsew signal tristate
flabel metal3 s 9517 8848 10317 8968 0 FreeSans 480 0 0 0 data_out[7]
port 10 nsew signal tristate
flabel metal2 s 5814 11661 5870 12461 0 FreeSans 224 90 0 0 in
port 11 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 rst
port 12 nsew signal input
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 rst_cap
port 13 nsew signal tristate
rlabel metal1 5152 9792 5152 9792 0 VGND
rlabel metal1 5152 9248 5152 9248 0 VPWR
rlabel metal1 4232 5338 4232 5338 0 _000_
rlabel via1 5009 3026 5009 3026 0 _001_
rlabel metal1 2330 2346 2330 2346 0 _002_
rlabel metal1 5244 4794 5244 4794 0 _003_
rlabel metal1 1886 8058 1886 8058 0 _004_
rlabel metal2 2990 8738 2990 8738 0 _005_
rlabel metal2 5750 8738 5750 8738 0 _006_
rlabel metal1 3910 6970 3910 6970 0 _007_
rlabel via1 1697 3026 1697 3026 0 _008_
rlabel via1 1697 4590 1697 4590 0 _009_
rlabel metal1 2484 5882 2484 5882 0 _010_
rlabel metal1 8372 3094 8372 3094 0 _011_
rlabel metal1 7912 3366 7912 3366 0 _012_
rlabel metal1 7774 2414 7774 2414 0 _013_
rlabel metal1 7866 5644 7866 5644 0 _014_
rlabel metal1 8234 4624 8234 4624 0 _015_
rlabel metal1 7636 4794 7636 4794 0 _016_
rlabel metal1 8556 6154 8556 6154 0 _017_
rlabel metal1 8694 6358 8694 6358 0 _018_
rlabel metal1 7820 7514 7820 7514 0 _019_
rlabel metal2 3910 5916 3910 5916 0 _020_
rlabel metal1 4600 2618 4600 2618 0 _021_
rlabel metal1 4140 3366 4140 3366 0 _022_
rlabel metal1 4554 3638 4554 3638 0 _023_
rlabel metal1 2944 2414 2944 2414 0 _024_
rlabel metal1 4048 6290 4048 6290 0 _025_
rlabel metal1 2645 7854 2645 7854 0 _026_
rlabel metal1 5336 4590 5336 4590 0 _027_
rlabel metal1 2300 7514 2300 7514 0 _028_
rlabel metal1 4002 7718 4002 7718 0 _029_
rlabel metal1 2622 7514 2622 7514 0 _030_
rlabel metal1 4094 7174 4094 7174 0 _031_
rlabel metal1 4278 6800 4278 6800 0 _032_
rlabel metal1 4646 7514 4646 7514 0 _033_
rlabel metal1 3588 6766 3588 6766 0 _034_
rlabel metal1 4554 6732 4554 6732 0 _035_
rlabel metal2 2990 4182 2990 4182 0 _036_
rlabel metal1 2162 5236 2162 5236 0 _037_
rlabel metal1 2162 3502 2162 3502 0 _038_
rlabel metal1 3312 5678 3312 5678 0 _039_
rlabel metal1 2346 5610 2346 5610 0 _040_
rlabel metal1 2254 5644 2254 5644 0 _041_
rlabel metal1 2622 5746 2622 5746 0 _042_
rlabel metal2 3818 7293 3818 7293 0 clk
rlabel metal2 5106 7174 5106 7174 0 clknet_0_clk
rlabel metal1 2254 2550 2254 2550 0 clknet_1_0__leaf_clk
rlabel metal1 3128 6766 3128 6766 0 clknet_1_1__leaf_clk
rlabel metal1 5842 6154 5842 6154 0 counter\[0\]
rlabel metal2 4646 3927 4646 3927 0 counter\[1\]
rlabel metal1 3726 2618 3726 2618 0 counter\[2\]
rlabel metal1 5290 4998 5290 4998 0 counter\[3\]
rlabel metal1 5842 7378 5842 7378 0 counter\[4\]
rlabel metal1 3036 7378 3036 7378 0 counter\[5\]
rlabel metal1 5244 7310 5244 7310 0 counter\[6\]
rlabel metal2 5842 8364 5842 8364 0 counter\[7\]
rlabel metal1 3128 4590 3128 4590 0 counter\[8\]
rlabel metal1 2990 5134 2990 5134 0 counter\[9\]
rlabel metal2 8694 3553 8694 3553 0 data_out[0]
rlabel metal1 8740 2618 8740 2618 0 data_out[1]
rlabel metal1 8924 4454 8924 4454 0 data_out[2]
rlabel metal2 8786 4913 8786 4913 0 data_out[3]
rlabel metal2 8694 6035 8694 6035 0 data_out[4]
rlabel metal1 8510 6834 8510 6834 0 data_out[5]
rlabel metal1 8924 7718 8924 7718 0 data_out[6]
rlabel metal2 8694 8993 8694 8993 0 data_out[7]
rlabel metal1 6210 9622 6210 9622 0 in
rlabel metal1 6026 9078 6026 9078 0 net1
rlabel metal1 8510 8976 8510 8976 0 net10
rlabel metal1 1656 6290 1656 6290 0 net11
rlabel metal1 2254 5168 2254 5168 0 net12
rlabel metal1 5106 2346 5106 2346 0 net13
rlabel metal1 5290 4454 5290 4454 0 net14
rlabel metal2 4370 6970 4370 6970 0 net15
rlabel metal2 2438 5916 2438 5916 0 net16
rlabel metal1 5060 2414 5060 2414 0 net17
rlabel metal1 3634 7990 3634 7990 0 net18
rlabel metal1 3082 8500 3082 8500 0 net19
rlabel metal1 4186 2380 4186 2380 0 net2
rlabel metal1 2530 7718 2530 7718 0 net20
rlabel metal1 8004 2618 8004 2618 0 net3
rlabel metal1 8142 2346 8142 2346 0 net4
rlabel metal1 8464 4590 8464 4590 0 net5
rlabel metal1 8464 5202 8464 5202 0 net6
rlabel metal1 8234 5678 8234 5678 0 net7
rlabel metal1 9016 6426 9016 6426 0 net8
rlabel metal1 8234 6834 8234 6834 0 net9
rlabel metal1 7866 2482 7866 2482 0 register_temp\[0\]
rlabel metal1 8050 3536 8050 3536 0 register_temp\[1\]
rlabel metal1 7314 4658 7314 4658 0 register_temp\[2\]
rlabel metal2 7774 4794 7774 4794 0 register_temp\[3\]
rlabel metal1 8280 6358 8280 6358 0 register_temp\[4\]
rlabel metal2 7774 6681 7774 6681 0 register_temp\[5\]
rlabel metal1 8050 7514 8050 7514 0 register_temp\[6\]
rlabel metal1 7544 8942 7544 8942 0 register_temp\[7\]
rlabel metal3 1050 7548 1050 7548 0 rst
rlabel metal3 751 6188 751 6188 0 rst_cap
<< properties >>
string FIXED_BBOX 0 0 10317 12461
<< end >>
