magic
tech sky130B
magscale 1 2
timestamp 1712303529
<< locali >>
rect 2148 3437 2303 3523
rect 2148 2894 2234 3437
rect 8772 1580 8876 1644
rect -1680 517 15526 552
rect -1680 466 2154 517
rect -1680 374 -914 466
rect -822 443 2154 466
rect 2228 443 15526 517
rect -822 374 15526 443
rect -1680 352 15526 374
rect -1694 -8 15808 192
<< viali >>
rect 2450 3588 2514 3652
rect 2630 3182 2666 3218
rect 2148 2788 2234 2874
rect 808 1880 872 1944
rect 7214 1580 7278 1644
rect 8708 1580 8772 1644
rect -914 374 -822 466
rect 2154 443 2228 517
<< metal1 >>
rect 2444 3658 2520 3664
rect 2444 3652 2456 3658
rect 2444 3588 2450 3652
rect 2444 3582 2456 3588
rect 2520 3582 2526 3658
rect 2444 3576 2520 3582
rect 2624 3226 2672 3230
rect 2616 3174 2622 3226
rect 2674 3174 2680 3226
rect 2624 3170 2672 3174
rect 2136 2874 2246 2880
rect 2136 2788 2148 2874
rect 2234 2788 2246 2874
rect 2136 2782 2246 2788
rect 802 1950 878 1956
rect 796 1874 802 1950
rect 866 1944 878 1950
rect 872 1880 878 1944
rect 866 1874 878 1880
rect 802 1868 878 1874
rect 2148 517 2234 2782
rect 7208 1650 7284 1656
rect 8702 1650 8778 1656
rect 7202 1586 7208 1650
rect 7284 1586 7290 1650
rect 7202 1580 7214 1586
rect 7278 1580 7290 1586
rect 7202 1574 7290 1580
rect 8696 1574 8702 1650
rect 8766 1644 8778 1650
rect 8772 1580 8778 1644
rect 8766 1574 8778 1580
rect 8702 1568 8778 1574
rect -920 472 -816 478
rect 2148 443 2154 517
rect 2228 443 2234 517
rect 2148 431 2234 443
rect -920 362 -816 368
<< via1 >>
rect 2456 3652 2520 3658
rect 2456 3588 2514 3652
rect 2514 3588 2520 3652
rect 2456 3582 2520 3588
rect 2622 3218 2674 3226
rect 2622 3182 2630 3218
rect 2630 3182 2666 3218
rect 2666 3182 2674 3218
rect 2622 3174 2674 3182
rect 802 1944 866 1950
rect 802 1880 808 1944
rect 808 1880 866 1944
rect 802 1874 866 1880
rect 7208 1644 7284 1650
rect 7208 1586 7214 1644
rect 7214 1586 7278 1644
rect 7278 1586 7284 1644
rect 8702 1644 8766 1650
rect 8702 1580 8708 1644
rect 8708 1580 8766 1644
rect 8702 1574 8766 1580
rect -920 466 -816 472
rect -920 374 -914 466
rect -914 374 -822 466
rect -822 374 -816 466
rect -920 368 -816 374
<< metal2 >>
rect 2456 3658 2520 3664
rect 2520 3588 2568 3652
rect 2632 3588 2641 3652
rect 2456 3576 2520 3582
rect 11788 3564 11852 3573
rect 11788 3491 11852 3500
rect 2622 3226 2674 3232
rect 2674 3182 2858 3218
rect 2622 3168 2674 3174
rect 802 1950 866 1956
rect 414 1880 802 1944
rect 802 1868 866 1874
rect 7008 1650 7072 1659
rect 8702 1650 8766 1656
rect 7072 1586 7208 1650
rect 7284 1586 7290 1650
rect 7008 1577 7072 1586
rect 8508 1580 8702 1644
rect 8702 1568 8766 1574
rect -926 368 -920 472
rect -816 368 -810 472
<< via2 >>
rect 2568 3588 2632 3652
rect 11788 3500 11852 3564
rect 7008 1586 7072 1650
rect -915 373 -821 467
<< metal3 >>
rect 2563 3652 2637 3657
rect 2563 3588 2568 3652
rect 2632 3588 2637 3652
rect 2563 3583 2637 3588
rect 2568 3092 2632 3583
rect 11788 3569 11852 4112
rect 11783 3564 11857 3569
rect 11783 3500 11788 3564
rect 11852 3500 11857 3564
rect 11783 3495 11857 3500
rect 7008 3092 7072 3098
rect 4222 3028 4228 3092
rect 4292 3028 4298 3092
rect 2568 3022 2632 3028
rect -920 471 -816 472
rect -925 369 -919 471
rect -817 369 -811 471
rect -920 368 -816 369
rect 2725 -108 2827 -103
rect 4228 -108 4292 3028
rect 7008 1655 7072 3028
rect 7003 1650 7077 1655
rect 7003 1586 7008 1650
rect 7072 1586 7077 1650
rect 7003 1581 7077 1586
rect 12373 -108 12475 -103
rect -4512 -109 17300 -108
rect -4517 -211 -4511 -109
rect -4409 -211 -2099 -109
rect -1997 -211 313 -109
rect 415 -211 2725 -109
rect 2827 -211 5137 -109
rect 5239 -211 7549 -109
rect 7651 -211 9961 -109
rect 10063 -211 12373 -109
rect 12475 -211 14785 -109
rect 14887 -211 17197 -109
rect 17299 -211 17305 -109
rect -4512 -212 17300 -211
rect 2725 -217 2827 -212
rect 12373 -217 12475 -212
rect -3338 -392 -3332 -288
rect -3228 -289 18492 -288
rect -3228 -391 -919 -289
rect -817 -391 1493 -289
rect 1595 -391 3905 -289
rect 4007 -391 6317 -289
rect 6419 -391 8729 -289
rect 8831 -391 11141 -289
rect 11243 -391 13553 -289
rect 13655 -391 15965 -289
rect 16067 -391 18377 -289
rect 18479 -391 18492 -289
rect -3228 -392 18492 -391
<< via3 >>
rect 2568 3028 2632 3092
rect 4228 3028 4292 3092
rect 7008 3028 7072 3092
rect -919 467 -817 471
rect -919 373 -915 467
rect -915 373 -821 467
rect -821 373 -817 467
rect -919 369 -817 373
rect -4511 -211 -4409 -109
rect -2099 -211 -1997 -109
rect 313 -211 415 -109
rect 2725 -211 2827 -109
rect 5137 -211 5239 -109
rect 7549 -211 7651 -109
rect 9961 -211 10063 -109
rect 12373 -211 12475 -109
rect 14785 -211 14887 -109
rect 17197 -211 17299 -109
rect -3332 -392 -3228 -288
rect -919 -391 -817 -289
rect 1493 -391 1595 -289
rect 3905 -391 4007 -289
rect 6317 -391 6419 -289
rect 8729 -391 8831 -289
rect 11141 -391 11243 -289
rect 13553 -391 13655 -289
rect 15965 -391 16067 -289
rect 18377 -391 18479 -289
<< metal4 >>
rect 2567 3092 2633 3093
rect 4227 3092 4293 3093
rect 7007 3092 7073 3093
rect 2548 3028 2568 3092
rect 2632 3028 4228 3092
rect 4292 3028 7008 3092
rect 7072 3028 7073 3092
rect 2567 3027 2633 3028
rect 4227 3027 4293 3028
rect 7007 3027 7073 3028
rect -920 471 -816 472
rect -920 369 -919 471
rect -817 369 -816 471
rect -4512 -109 -4408 -108
rect -4512 -211 -4511 -109
rect -4409 -211 -4408 -109
rect -4512 -512 -4408 -211
rect -2100 -109 -1996 -108
rect -2100 -211 -2099 -109
rect -1997 -211 -1996 -109
rect -3333 -288 -3227 -287
rect -3333 -392 -3332 -288
rect -3228 -392 -3227 -288
rect -3333 -393 -3227 -392
rect -3332 -512 -3228 -393
rect -2100 -512 -1996 -211
rect -920 -289 -816 369
rect -920 -391 -919 -289
rect -817 -391 -816 -289
rect -920 -512 -816 -391
rect 312 -109 416 -108
rect 312 -211 313 -109
rect 415 -211 416 -109
rect 312 -504 416 -211
rect 2724 -109 2828 -108
rect 2724 -211 2725 -109
rect 2827 -211 2828 -109
rect 1492 -289 1596 -288
rect 1492 -391 1493 -289
rect 1595 -391 1596 -289
rect 1492 -512 1596 -391
rect 2724 -504 2828 -211
rect 5136 -109 5240 -108
rect 5136 -211 5137 -109
rect 5239 -211 5240 -109
rect 3904 -289 4008 -288
rect 3904 -391 3905 -289
rect 4007 -391 4008 -289
rect 3904 -504 4008 -391
rect 5136 -512 5240 -211
rect 7548 -109 7652 -108
rect 7548 -211 7549 -109
rect 7651 -211 7652 -109
rect 6316 -289 6420 -288
rect 6316 -391 6317 -289
rect 6419 -391 6420 -289
rect 6316 -504 6420 -391
rect 7548 -504 7652 -211
rect 9960 -109 10064 -108
rect 9960 -211 9961 -109
rect 10063 -211 10064 -109
rect 8728 -289 8832 -288
rect 8728 -391 8729 -289
rect 8831 -391 8832 -289
rect 8728 -512 8832 -391
rect 9960 -504 10064 -211
rect 12372 -109 12476 -108
rect 12372 -211 12373 -109
rect 12475 -211 12476 -109
rect 11140 -289 11244 -288
rect 11140 -391 11141 -289
rect 11243 -391 11244 -289
rect 11140 -532 11244 -391
rect 12372 -504 12476 -211
rect 14784 -109 14888 -108
rect 14784 -211 14785 -109
rect 14887 -211 14888 -109
rect 13552 -289 13656 -288
rect 13552 -391 13553 -289
rect 13655 -391 13656 -289
rect 13552 -504 13656 -391
rect 14784 -504 14888 -211
rect 17196 -109 17300 -108
rect 17196 -211 17197 -109
rect 17299 -211 17300 -109
rect 15964 -289 16068 -288
rect 15964 -391 15965 -289
rect 16067 -391 16068 -289
rect 15964 -512 16068 -391
rect 17196 -512 17300 -211
rect 18376 -289 18480 -288
rect 18376 -391 18377 -289
rect 18479 -391 18480 -289
rect 18376 -532 18480 -391
use CM_OTA_NCH  CM_OTA_NCH_0
timestamp 1712302962
transform 1 0 7606 0 1 1092
box -7620 -1100 8200 5936
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 2184 -1 0 4228
box -184 -124 1528 728
use sky130_fd_pr__cap_mim_m3_1_TWL4V4  sky130_fd_pr__cap_mim_m3_1_TWL4V4_0
timestamp 1711374513
transform 1 0 6540 0 1 -5900
box -11940 -5500 11940 5500
<< labels >>
flabel metal2 2674 3182 2858 3218 0 FreeSans 800 0 0 0 RST
port 1 nsew
flabel metal3 11788 3564 11852 4112 0 FreeSans 800 0 0 0 OUT
port 2 nsew
flabel metal4 2632 3028 7008 3092 0 FreeSans 800 0 0 0 I_IN
port 3 nsew
flabel metal2 8508 1580 8702 1644 0 FreeSans 800 0 0 0 VREF_I
port 4 nsew
flabel locali -1680 -8 4480 192 0 FreeSans 800 0 0 0 VDD
port 5 nsew
flabel locali -1680 352 12286 552 0 FreeSans 800 0 0 0 VSS
port 6 nsew
flabel metal2 414 1880 802 1944 0 FreeSans 800 0 0 0 IBIAS
port 7 nsew
<< end >>
