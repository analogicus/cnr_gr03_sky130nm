magic
tech sky130B
magscale 1 2
timestamp 1712848679
<< locali >>
rect 2295 5039 2399 5102
rect 2295 5033 2381 5039
rect -5512 3378 -4704 3598
rect 252 2786 324 3186
rect 956 2750 1020 3252
rect 2596 2740 2660 4732
rect 4023 3906 4658 3992
rect 4023 3835 4109 3906
rect 3900 3534 3964 3538
rect 3900 3482 3914 3534
rect 3900 3384 3964 3482
rect 5631 3434 6054 3506
rect 3900 3320 4380 3384
rect 3612 2780 3684 3186
rect 4316 2736 4380 3250
rect 2180 2644 2656 2708
rect 2180 2522 2244 2644
rect 252 1770 324 2166
rect 956 1722 1020 2230
rect 3612 1794 3684 2262
rect 6265 2243 6409 2329
rect 4316 2032 4380 2230
rect 4316 1722 4380 1968
rect 6323 1694 6409 2243
rect 2180 1566 2662 1630
rect 2180 1502 2244 1566
rect 2180 1434 2244 1438
rect 956 1204 1020 1210
rect 956 1152 966 1204
rect 1018 1152 1020 1204
rect 252 730 324 1146
rect 956 698 1020 1152
rect 2305 1074 2391 1137
rect 2305 988 2887 1074
rect 3612 774 3684 1276
rect 4316 712 4380 1218
rect 5108 653 5253 739
rect 5108 109 5194 653
rect -5528 -579 7300 -374
rect -5528 -653 2893 -579
rect 2967 -653 7300 -579
rect -5528 -792 7300 -653
rect -5536 -1181 7292 -1000
rect -5536 -1255 4635 -1181
rect 4709 -1212 6329 -1181
rect 4709 -1255 5328 -1212
rect -5536 -1264 5328 -1255
rect 5380 -1255 6329 -1212
rect 6403 -1255 7292 -1181
rect 5380 -1264 7292 -1255
rect -5536 -1418 7292 -1264
<< viali >>
rect 2232 4824 2284 4876
rect 1944 4610 1996 4662
rect -1004 3444 -952 3496
rect 252 3438 316 3502
rect 540 3474 604 3538
rect 3914 3482 3966 3534
rect 5478 2772 5542 2836
rect 6094 2772 6158 2836
rect 540 2456 604 2520
rect 2180 2458 2244 2522
rect 3910 2464 3962 2516
rect 2186 2108 2238 2160
rect 4316 1968 4380 2032
rect 5436 1974 5488 2026
rect 6030 1974 6082 2026
rect 6323 1588 6409 1674
rect 540 1432 604 1496
rect 2180 1438 2244 1502
rect 3900 1438 3964 1502
rect 966 1152 1018 1204
rect 2596 1146 2660 1210
rect 2887 988 2973 1074
rect 6136 760 6188 812
rect 546 428 598 480
rect 3900 414 3964 478
rect 5322 392 5386 456
rect 4629 -32 4715 54
rect 2893 -653 2967 -579
rect 4635 -1255 4709 -1181
rect 5328 -1264 5380 -1212
rect 6329 -1255 6403 -1181
<< metal1 >>
rect 2226 4876 2290 4888
rect 2226 4824 2232 4876
rect 2284 4824 2290 4876
rect 1938 4662 2002 4674
rect 1938 4610 1944 4662
rect 1996 4610 2002 4662
rect 528 3538 616 3544
rect 246 3508 322 3514
rect -1010 3502 -946 3508
rect -1010 3432 -946 3438
rect 240 3432 246 3508
rect 310 3502 322 3508
rect 316 3438 322 3502
rect 528 3474 540 3538
rect 604 3474 616 3538
rect 528 3468 616 3474
rect 310 3432 322 3438
rect 246 3426 322 3432
rect 540 3326 604 3468
rect 1938 3326 2002 4610
rect 2226 3540 2290 4824
rect 2226 3470 2290 3476
rect 3908 3540 3972 3546
rect 3908 3470 3972 3476
rect 534 3262 540 3326
rect 604 3262 610 3326
rect 540 2526 604 3262
rect 1938 3256 2002 3262
rect 5472 2842 5548 2848
rect 5472 2836 5484 2842
rect 5472 2772 5478 2836
rect 5472 2766 5484 2772
rect 5548 2766 5554 2842
rect 6082 2836 6170 2842
rect 5754 2772 5760 2836
rect 5824 2772 5830 2836
rect 6082 2772 6094 2836
rect 6158 2772 6170 2836
rect 5472 2760 5548 2766
rect 2174 2528 2250 2534
rect 534 2520 610 2526
rect 534 2456 540 2520
rect 604 2456 610 2520
rect 534 2450 610 2456
rect 2174 2522 2186 2528
rect 2174 2458 2180 2522
rect 2174 2452 2186 2458
rect 2250 2452 2256 2528
rect 3904 2522 3968 2528
rect 3904 2452 3968 2458
rect 540 1502 604 2450
rect 2174 2446 2250 2452
rect 2180 2160 2244 2172
rect 2180 2108 2186 2160
rect 2238 2108 2244 2160
rect 2180 2008 2244 2108
rect 2742 2106 2748 2170
rect 2812 2106 2818 2170
rect 2748 2008 2812 2106
rect 4310 2038 4386 2044
rect 4310 2032 4322 2038
rect 2742 1944 2748 2008
rect 2812 1944 2818 2008
rect 4310 1968 4316 2032
rect 4310 1962 4322 1968
rect 4386 1962 4392 2038
rect 5430 2032 5494 2038
rect 5760 2032 5824 2772
rect 6082 2766 6170 2772
rect 6094 2170 6158 2766
rect 6088 2106 6094 2170
rect 6158 2106 6164 2170
rect 6024 2032 6088 2038
rect 5754 1968 5760 2032
rect 5824 1968 5830 2032
rect 5430 1962 5494 1968
rect 4310 1956 4386 1962
rect 2180 1508 2244 1944
rect 2168 1502 2256 1508
rect 534 1496 610 1502
rect 534 1432 540 1496
rect 604 1432 610 1496
rect 2168 1438 2180 1502
rect 2244 1438 2256 1502
rect 2168 1432 2256 1438
rect 3888 1502 3976 1508
rect 3888 1438 3900 1502
rect 3964 1438 3976 1502
rect 3888 1432 3976 1438
rect 534 1426 610 1432
rect 540 480 604 1426
rect 3900 1240 3964 1432
rect 2590 1216 2666 1222
rect 960 1210 1024 1216
rect 960 1140 1024 1146
rect 2584 1140 2590 1216
rect 2654 1210 2666 1216
rect 2660 1146 2666 1210
rect 2654 1140 2666 1146
rect 2590 1134 2666 1140
rect 5760 1102 5824 1968
rect 6024 1962 6088 1968
rect 6311 1674 6421 1680
rect 6311 1588 6323 1674
rect 6409 1588 6421 1674
rect 6311 1582 6421 1588
rect 2875 1074 2985 1080
rect 2875 988 2887 1074
rect 2973 988 2985 1074
rect 5754 1038 5760 1102
rect 5824 1038 5830 1102
rect 6124 1038 6130 1102
rect 6194 1038 6200 1102
rect 2875 982 2985 988
rect 540 428 546 480
rect 598 428 604 480
rect 540 416 604 428
rect 2887 -579 2973 982
rect 6130 812 6194 1038
rect 6130 760 6136 812
rect 6188 760 6194 812
rect 6130 748 6194 760
rect 3888 478 3976 484
rect 3888 414 3900 478
rect 3964 414 3976 478
rect 3888 408 3976 414
rect 5310 456 5398 462
rect 3900 220 3964 408
rect 5310 392 5322 456
rect 5386 392 5398 456
rect 5310 386 5398 392
rect 4617 54 4727 60
rect 4617 -32 4629 54
rect 4715 -32 4727 54
rect 4617 -38 4727 -32
rect 2887 -653 2893 -579
rect 2967 -653 2973 -579
rect 2887 -665 2973 -653
rect 4629 -1181 4715 -38
rect 4629 -1255 4635 -1181
rect 4709 -1255 4715 -1181
rect 4629 -1267 4715 -1255
rect 5322 -1212 5386 386
rect 5322 -1264 5328 -1212
rect 5380 -1264 5386 -1212
rect 5322 -1276 5386 -1264
rect 6323 -1181 6409 1582
rect 6323 -1255 6329 -1181
rect 6403 -1255 6409 -1181
rect 6323 -1267 6409 -1255
<< via1 >>
rect -1010 3496 -946 3502
rect -1010 3444 -1004 3496
rect -1004 3444 -952 3496
rect -952 3444 -946 3496
rect -1010 3438 -946 3444
rect 246 3502 310 3508
rect 246 3438 252 3502
rect 252 3438 310 3502
rect 246 3432 310 3438
rect 2226 3476 2290 3540
rect 3908 3534 3972 3540
rect 3908 3482 3914 3534
rect 3914 3482 3966 3534
rect 3966 3482 3972 3534
rect 3908 3476 3972 3482
rect 540 3262 604 3326
rect 1938 3262 2002 3326
rect 5484 2836 5548 2842
rect 5484 2772 5542 2836
rect 5542 2772 5548 2836
rect 5484 2766 5548 2772
rect 5760 2772 5824 2836
rect 2186 2522 2250 2528
rect 2186 2458 2244 2522
rect 2244 2458 2250 2522
rect 2186 2452 2250 2458
rect 3904 2516 3968 2522
rect 3904 2464 3910 2516
rect 3910 2464 3962 2516
rect 3962 2464 3968 2516
rect 3904 2458 3968 2464
rect 2748 2106 2812 2170
rect 4322 2032 4386 2038
rect 2180 1944 2244 2008
rect 2748 1944 2812 2008
rect 4322 1968 4380 2032
rect 4380 1968 4386 2032
rect 4322 1962 4386 1968
rect 6094 2106 6158 2170
rect 5430 2026 5494 2032
rect 5430 1974 5436 2026
rect 5436 1974 5488 2026
rect 5488 1974 5494 2026
rect 5430 1968 5494 1974
rect 5760 1968 5824 2032
rect 6024 2026 6088 2032
rect 6024 1974 6030 2026
rect 6030 1974 6082 2026
rect 6082 1974 6088 2026
rect 6024 1968 6088 1974
rect 960 1204 1024 1210
rect 960 1152 966 1204
rect 966 1152 1018 1204
rect 1018 1152 1024 1204
rect 960 1146 1024 1152
rect 2590 1210 2654 1216
rect 2590 1146 2596 1210
rect 2596 1146 2654 1210
rect 2590 1140 2654 1146
rect 5760 1038 5824 1102
rect 6130 1038 6194 1102
<< metal2 >>
rect 246 3508 310 3514
rect -1016 3438 -1010 3502
rect -946 3438 246 3502
rect 2220 3476 2226 3540
rect 2290 3476 3908 3540
rect 3972 3476 3978 3540
rect 246 3426 310 3432
rect 540 3326 604 3332
rect 604 3262 1938 3326
rect 2002 3262 2008 3326
rect 540 3256 604 3262
rect 5484 2842 5548 2848
rect 5760 2836 5824 2842
rect 5548 2772 5760 2836
rect 5760 2766 5824 2772
rect 5484 2760 5548 2766
rect 2186 2528 2250 2534
rect 2250 2458 3904 2522
rect 3968 2458 3974 2522
rect 2186 2446 2250 2452
rect 2748 2170 2812 2176
rect 6094 2170 6158 2176
rect 2812 2106 6094 2170
rect 2748 2100 2812 2106
rect 6094 2100 6158 2106
rect 4322 2038 4386 2044
rect 2748 2008 2812 2014
rect 2174 1944 2180 2008
rect 2244 1944 2748 2008
rect 5760 2032 5824 2038
rect 4386 1968 5430 2032
rect 5494 1968 5500 2032
rect 5824 1968 6024 2032
rect 6088 1968 6094 2032
rect 5760 1962 5824 1968
rect 4322 1956 4386 1962
rect 2748 1938 2812 1944
rect 2590 1216 2654 1222
rect 954 1146 960 1210
rect 1024 1146 2590 1210
rect 2590 1134 2654 1140
rect 5760 1102 5824 1108
rect 6130 1102 6194 1108
rect 5824 1038 6130 1102
rect 5760 1032 5824 1038
rect 6130 1032 6194 1038
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 5144 -1 0 1256
box -184 -124 1336 2168
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 1606 0 1 4548
box -184 -124 1528 728
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 1604 0 1 1024
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_2
timestamp 1695852000
transform 1 0 1604 0 1 2044
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_3
timestamp 1695852000
transform 1 0 -36 0 1 4
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_4
timestamp 1695852000
transform 1 0 -36 0 1 3064
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_5
timestamp 1695852000
transform 1 0 -36 0 1 2044
box -184 -124 1528 1016
use CNRATR_NCH_4C4F0  CNRATR_NCH_4C4F0_6
timestamp 1695852000
transform 1 0 -36 0 1 1024
box -184 -124 1528 1016
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 1 0 3324 0 1 4
box -184 -124 1528 1016
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_1
timestamp 1695852000
transform 1 0 3324 0 1 3064
box -184 -124 1528 1016
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_2
timestamp 1695852000
transform 1 0 3324 0 1 2044
box -184 -124 1528 1016
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_3
timestamp 1695852000
transform 1 0 3324 0 1 1024
box -184 -124 1528 1016
use CNRATR_PCH_12C1F2  CNRATR_PCH_12C1F2_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 5884 -1 0 3796
box -184 -124 2296 613
use CNRATR_PCH_12C1F2  CNRATR_PCH_12C1F2_1
timestamp 1695852000
transform 0 1 5264 -1 0 3796
box -184 -124 2296 613
use SUNTR_RPPO8  SUNTR_RPPO8_0 ~/aicex/ip/cnr_gr03_sky130nm/design/SUN_TR_SKY130NM
timestamp 1712819652
transform 1 0 -5540 0 1 -60
box 0 0 5264 4236
<< labels >>
flabel locali -5528 -792 7300 -374 0 FreeSans 800 0 0 0 VSS
port 2 nsew
flabel locali -5536 -1418 7292 -1000 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel metal1 3900 1240 3964 1438 0 FreeSans 800 0 0 0 IBIAS1_2u
port 3 nsew
flabel metal1 3900 220 3964 414 0 FreeSans 800 0 0 0 IBIAS2_2u
port 4 nsew
<< end >>
