magic
tech sky130B
magscale 1 2
timestamp 1710170680
<< locali >>
rect -150 5350 40 5400
rect 1300 5350 1490 5400
rect 2780 5350 2970 5400
rect -1550 4504 -1420 4544
rect -1550 3960 -1510 4504
rect 4241 4505 4389 4544
rect -230 4260 100 4310
rect 2710 4260 3060 4310
rect 4350 3991 4389 4505
rect 4960 3930 5010 4240
rect 5660 3980 5720 4180
rect 6560 3930 6610 4230
rect 7260 3980 7320 4180
rect 4960 3330 5010 3640
rect 5660 3380 5720 3580
rect 6560 3330 6610 3640
rect 7260 3380 7320 3580
rect -5666 2828 -5434 2900
rect -4786 2824 -4544 2896
rect -77 2660 -31 2871
rect 4960 2730 5010 3040
rect 5660 2780 5720 2980
rect 6560 2730 6610 3040
rect 7260 2780 7320 2980
rect -6472 2367 -6317 2453
rect -6472 1854 -6386 2367
rect -6020 2130 -5956 2502
rect -5738 2132 -5368 2196
rect -3680 2140 -3620 2434
rect -2753 2367 -2596 2453
rect -2682 1854 -2596 2367
rect 1040 2290 1330 2340
rect 1630 2290 1920 2340
rect 2220 2290 2510 2340
rect 4960 2130 5010 2440
rect 5660 2180 5720 2380
rect 6560 2130 6610 2440
rect 7260 2180 7320 2380
rect -500 1960 -190 2010
rect 4674 1648 4727 1734
rect 6274 1648 6577 1734
rect -5590 1068 -5354 1140
rect -4130 1068 -3894 1140
rect -2670 946 -2598 1066
rect 5600 1064 5846 1136
rect -2670 894 -2294 946
rect -2666 874 -2294 894
rect 970 876 1174 948
rect -6232 788 -5928 852
rect -6972 617 -6817 703
rect -6972 94 -6886 617
rect -5992 388 -5928 788
rect -494 659 -444 660
rect -494 628 -431 659
rect -489 569 -431 628
rect -319 569 -261 679
rect 2467 607 2628 693
rect -489 511 -261 569
rect -5672 372 -5258 436
rect -4202 372 -3798 436
rect -5518 0 -5426 80
rect -6070 -540 -4980 0
rect -2590 -10 -2400 180
rect -408 91 -350 511
rect 2542 180 2628 607
rect 2745 619 2895 669
rect 2745 180 2795 619
rect 7063 617 7207 671
rect 5518 372 5912 436
rect 2542 94 2795 180
rect 7153 123 7207 617
rect 2600 55 2795 94
rect -120 -540 960 10
rect 2600 -10 2790 55
rect 6010 -540 7100 0
rect -7100 -583 8200 -540
rect -7100 -593 6583 -583
rect -7100 -666 4734 -593
rect 4807 -657 6583 -593
rect 6657 -657 8200 -583
rect 4807 -666 8200 -657
rect -7100 -740 8200 -666
rect -7100 -877 8200 -850
rect -7100 -906 559 -877
rect -7100 -913 -1543 -906
rect -7100 -987 -6466 -913
rect -6392 -918 -1543 -913
rect -6392 -982 -2670 -918
rect -2606 -974 -1543 -918
rect -1475 -942 559 -906
rect 624 -883 8200 -877
rect 624 -942 2914 -883
rect -1475 -957 2914 -942
rect 2988 -904 8200 -883
rect 2988 -957 4309 -904
rect -1475 -974 4309 -957
rect -2606 -976 4309 -974
rect 4381 -976 8200 -904
rect -2606 -982 8200 -976
rect -6392 -987 8200 -982
rect -7100 -1050 8200 -987
<< viali >>
rect -814 4490 -746 4558
rect 657 4501 704 4548
rect 2110 4494 2171 4555
rect 3603 4507 3637 4541
rect 2355 4255 2404 4304
rect 5368 4350 5432 4384
rect 6968 4350 7032 4387
rect -1552 3868 -1466 3954
rect 4302 3868 4388 3954
rect 5383 3763 5417 3797
rect 6984 3774 7018 3808
rect 5384 3164 5418 3198
rect 6968 3158 7032 3194
rect -808 3052 -752 3108
rect 136 3036 185 3085
rect 663 2993 698 3028
rect 1656 3016 1728 3050
rect 2414 3004 2448 3038
rect -90 2900 -29 2961
rect 860 2710 900 2750
rect 2030 2698 2094 2762
rect 1093 2537 1127 2571
rect 1463 2537 1497 2571
rect 1833 2533 1867 2567
rect 2640 2534 2680 2574
rect 5384 2563 5418 2597
rect 6984 2563 7018 2597
rect -5141 2408 -5098 2451
rect -3305 2134 -3254 2185
rect -689 2195 -630 2254
rect -90 2194 -30 2254
rect 548 1898 634 1975
rect 2908 1898 2994 1984
rect 5384 1963 5418 1997
rect 6984 1963 7018 1997
rect -6472 1748 -6386 1834
rect -2682 1748 -2596 1834
rect 5648 1734 5720 1806
rect 7248 1734 7320 1806
rect 4727 1648 4813 1734
rect 6577 1648 6663 1734
rect -4768 932 -4713 987
rect -3312 964 -3248 1028
rect 3470 960 3530 1020
rect 1174 876 1246 948
rect 4960 940 5020 1000
rect 6420 950 6480 1010
rect -1429 775 -1371 833
rect 330 774 390 834
rect 1831 775 1889 833
rect 4734 -666 4807 -593
rect 6583 -657 6657 -583
rect -6466 -987 -6392 -913
rect -2670 -982 -2606 -918
rect -1543 -974 -1475 -906
rect 559 -942 624 -877
rect 2914 -957 2988 -883
rect 4309 -976 4381 -904
<< metal1 >>
rect -826 4558 -734 4564
rect -826 4490 -814 4558
rect -746 4490 -734 4558
rect 2098 4555 2183 4561
rect 645 4548 716 4554
rect 645 4501 657 4548
rect 704 4501 716 4548
rect 645 4495 716 4501
rect -826 4484 -734 4490
rect -1564 3954 -1454 3960
rect -1564 3868 -1552 3954
rect -1466 3868 -1454 3954
rect -1564 3862 -1454 3868
rect -6028 2328 -5971 2468
rect -6028 2265 -5971 2271
rect -5147 2451 -5092 2463
rect -5147 2408 -5141 2451
rect -5098 2408 -5092 2451
rect -5147 2027 -5092 2408
rect -4774 2271 -4768 2328
rect -4711 2271 -4705 2328
rect -5147 1966 -5092 1972
rect -6484 1834 -6374 1840
rect -6484 1748 -6472 1834
rect -6386 1748 -6374 1834
rect -6484 1742 -6374 1748
rect -6472 -913 -6386 1742
rect -4768 993 -4711 2271
rect -3311 2185 -3248 2197
rect -3311 2134 -3305 2185
rect -3254 2134 -3248 2185
rect -3311 1034 -3248 2134
rect -2694 1834 -2584 1840
rect -2694 1748 -2682 1834
rect -2596 1748 -2584 1834
rect -2694 1742 -2584 1748
rect -3324 1028 -3236 1034
rect -4780 987 -4701 993
rect -4780 932 -4768 987
rect -4713 932 -4701 987
rect -3324 964 -3312 1028
rect -3248 964 -3236 1028
rect -3324 958 -3236 964
rect -4780 926 -4701 932
rect -2677 -208 -2600 1742
rect -1550 1719 -1468 3862
rect -814 3108 -746 4484
rect 124 3730 130 3791
rect 191 3730 197 3791
rect -814 3052 -808 3108
rect -752 3052 -746 3108
rect -814 3040 -746 3052
rect 130 3085 191 3730
rect 130 3036 136 3085
rect 185 3036 191 3085
rect 130 3024 191 3036
rect 269 3650 330 3656
rect -96 2967 -23 2973
rect -96 2961 -84 2967
rect -96 2900 -90 2961
rect -96 2894 -84 2900
rect -23 2894 -17 2967
rect 269 2961 330 3589
rect 657 3028 704 4495
rect 2098 4494 2110 4555
rect 2171 4494 2183 4555
rect 3591 4541 3649 4547
rect 3591 4507 3603 4541
rect 3637 4507 3649 4541
rect 3591 4501 3649 4507
rect 2098 4488 2183 4494
rect 2110 3791 2171 4488
rect 2110 3724 2171 3730
rect 2349 4304 2410 4316
rect 2349 4255 2355 4304
rect 2404 4255 2410 4304
rect 2349 3650 2410 4255
rect 2343 3589 2349 3650
rect 2410 3589 2416 3650
rect 3604 3363 3637 4501
rect 5356 4384 5444 4390
rect 5356 4350 5368 4384
rect 5432 4350 5444 4384
rect 5356 4344 5444 4350
rect 6956 4387 7044 4393
rect 6956 4350 6968 4387
rect 7032 4350 7044 4387
rect 6956 4344 7044 4350
rect 4290 3954 4400 3960
rect 4290 3868 4302 3954
rect 4388 3868 4400 3954
rect 4290 3862 4400 3868
rect 3595 3357 3647 3363
rect 2398 3305 2404 3357
rect 2456 3305 2462 3357
rect 1924 3236 1976 3242
rect 1924 3178 1976 3184
rect 1661 3104 1667 3156
rect 1719 3104 1725 3156
rect 1676 3056 1709 3104
rect 657 2993 663 3028
rect 698 2993 704 3028
rect 1644 3050 1740 3056
rect 1644 3016 1656 3050
rect 1728 3016 1740 3050
rect 1644 3010 1740 3016
rect 657 2981 704 2993
rect 269 2894 330 2900
rect -96 2888 -23 2894
rect 854 2756 906 2762
rect 1931 2756 1969 3178
rect 2414 3163 2446 3305
rect 3595 3299 3647 3305
rect 3754 3346 3806 3352
rect 3754 3288 3806 3294
rect 3761 3236 3799 3288
rect 3748 3184 3754 3236
rect 3806 3184 3812 3236
rect 2404 3157 2456 3163
rect 2404 3099 2456 3105
rect 2414 3050 2447 3099
rect 2408 3038 2454 3050
rect 3958 3044 3964 3096
rect 4016 3044 4022 3096
rect 2408 3004 2414 3038
rect 2448 3004 2454 3038
rect 2408 2992 2454 3004
rect 2024 2768 2100 2774
rect 1918 2704 1924 2756
rect 1976 2704 1982 2756
rect 854 2698 906 2704
rect 2018 2692 2024 2768
rect 2088 2762 2100 2768
rect 2094 2698 2100 2762
rect 2088 2692 2100 2698
rect 2024 2686 2100 2692
rect 1457 2580 1503 2583
rect 2634 2580 2686 2586
rect 1081 2571 1139 2577
rect 1081 2537 1093 2571
rect 1127 2537 1139 2571
rect 1081 2531 1139 2537
rect 1094 2452 1126 2531
rect 1448 2528 1454 2580
rect 1506 2528 1512 2580
rect 1827 2567 1873 2579
rect 1827 2533 1833 2567
rect 1867 2533 1873 2567
rect 1457 2525 1503 2528
rect 1827 2521 1873 2533
rect 2498 2528 2504 2580
rect 2556 2528 2562 2580
rect 1084 2446 1136 2452
rect 1834 2446 1866 2521
rect 2514 2456 2546 2528
rect 2634 2522 2686 2528
rect 3974 2462 4006 3044
rect 3964 2456 4016 2462
rect 1818 2394 1824 2446
rect 1876 2394 1882 2446
rect 2498 2404 2504 2456
rect 2556 2404 2562 2456
rect 3964 2398 4016 2404
rect 1084 2388 1136 2394
rect -701 2254 -618 2260
rect -701 2195 -689 2254
rect -630 2195 -618 2254
rect -701 2189 -618 2195
rect -102 2254 -18 2260
rect -102 2194 -90 2254
rect -30 2194 -18 2254
rect -1433 1972 -1427 2027
rect -1372 1972 -1366 2027
rect -6472 -987 -6466 -913
rect -6392 -987 -6386 -913
rect -6472 -999 -6386 -987
rect -2676 -918 -2600 -208
rect -1549 -900 -1469 1719
rect -1427 845 -1372 1972
rect -688 1400 -629 2189
rect -102 2188 -18 2194
rect -90 1490 -30 2188
rect 2896 1984 3006 1990
rect 536 1975 646 1981
rect 536 1898 548 1975
rect 634 1898 646 1975
rect 536 1892 646 1898
rect 2896 1898 2908 1984
rect 2994 1898 3006 1984
rect 2896 1892 3006 1898
rect -90 1424 -30 1430
rect -688 1335 -629 1341
rect 329 1400 392 1410
rect 329 1341 330 1400
rect 389 1341 392 1400
rect 329 1053 392 1341
rect -1435 833 -1365 845
rect 327 840 393 1053
rect -1435 775 -1429 833
rect -1371 775 -1365 833
rect -1435 763 -1365 775
rect 318 834 402 840
rect 318 774 330 834
rect 390 774 402 834
rect 318 768 402 774
rect 553 -877 630 1892
rect 1830 1490 1890 1496
rect 1830 1340 1890 1430
rect 1174 1276 1246 1282
rect 1174 954 1246 1204
rect 1162 948 1258 954
rect 1162 876 1174 948
rect 1246 876 1258 948
rect 1162 870 1258 876
rect 1831 839 1889 1340
rect 1819 833 1901 839
rect 1819 775 1831 833
rect 1889 775 1901 833
rect 1819 769 1901 775
rect -2676 -982 -2670 -918
rect -2606 -982 -2600 -918
rect -1555 -906 -1463 -900
rect -1555 -974 -1543 -906
rect -1475 -974 -1463 -906
rect 553 -942 559 -877
rect 624 -942 630 -877
rect 553 -954 630 -942
rect 2908 -883 2994 1892
rect 3458 1204 3464 1276
rect 3536 1204 3542 1276
rect 3464 1026 3536 1204
rect 3458 1020 3542 1026
rect 3458 960 3470 1020
rect 3530 960 3542 1020
rect 3458 954 3542 960
rect 2908 -957 2914 -883
rect 2988 -957 2994 -883
rect 2908 -969 2994 -957
rect 4303 -904 4387 3862
rect 5386 3809 5414 4344
rect 6985 3820 7016 4344
rect 5377 3797 5423 3809
rect 5377 3763 5383 3797
rect 5417 3763 5423 3797
rect 5377 3751 5423 3763
rect 6978 3808 7024 3820
rect 6978 3774 6984 3808
rect 7018 3774 7024 3808
rect 6978 3762 7024 3774
rect 5384 3210 5417 3751
rect 6984 3346 7018 3762
rect 6968 3294 6974 3346
rect 7026 3294 7032 3346
rect 5378 3198 5424 3210
rect 6984 3200 7018 3294
rect 5378 3164 5384 3198
rect 5418 3164 5424 3198
rect 5378 3152 5424 3164
rect 6956 3194 7044 3200
rect 6956 3158 6968 3194
rect 7032 3158 7044 3194
rect 6956 3152 7044 3158
rect 5384 3102 5418 3152
rect 5374 3096 5426 3102
rect 5374 3038 5426 3044
rect 5384 2609 5418 3038
rect 6984 2609 7018 3152
rect 5378 2597 5424 2609
rect 5378 2563 5384 2597
rect 5418 2563 5424 2597
rect 5378 2551 5424 2563
rect 6978 2597 7024 2609
rect 6978 2563 6984 2597
rect 7018 2563 7024 2597
rect 6978 2551 7024 2563
rect 5384 2009 5418 2551
rect 6984 2009 7018 2551
rect 5378 1997 5424 2009
rect 5378 1963 5384 1997
rect 5418 1963 5424 1997
rect 5378 1951 5424 1963
rect 6978 1997 7024 2009
rect 6978 1963 6984 1997
rect 7018 1963 7024 1997
rect 6978 1951 7024 1963
rect 5636 1806 5732 1812
rect 4721 1734 4819 1746
rect 4721 1648 4727 1734
rect 4813 1648 4819 1734
rect 5636 1734 5648 1806
rect 5720 1734 5732 1806
rect 7236 1806 7332 1812
rect 5636 1728 5732 1734
rect 6571 1734 6669 1746
rect 4721 1636 4819 1648
rect 4728 -593 4813 1636
rect 4954 1276 5026 1282
rect 4954 1000 5026 1204
rect 5648 1276 5720 1728
rect 6571 1648 6577 1734
rect 6663 1648 6669 1734
rect 7236 1734 7248 1806
rect 7320 1734 7332 1806
rect 7236 1728 7332 1734
rect 6571 1636 6669 1648
rect 6408 1204 6414 1276
rect 6486 1204 6492 1276
rect 5648 1198 5720 1204
rect 4954 940 4960 1000
rect 5020 940 5026 1000
rect 4954 928 5026 940
rect 6414 1010 6486 1204
rect 6414 950 6420 1010
rect 6480 950 6486 1010
rect 6414 938 6486 950
rect 4728 -666 4734 -593
rect 4807 -666 4813 -593
rect 4728 -678 4813 -666
rect 6577 -583 6663 1636
rect 7248 1276 7320 1728
rect 7248 1198 7320 1204
rect 6577 -657 6583 -583
rect 6657 -657 6663 -583
rect 6577 -669 6663 -657
rect -1555 -980 -1463 -974
rect 4303 -976 4309 -904
rect 4381 -976 4387 -904
rect -2676 -994 -2600 -982
rect 4303 -988 4387 -976
<< via1 >>
rect -6028 2271 -5971 2328
rect -4768 2271 -4711 2328
rect -5147 1972 -5092 2027
rect 130 3730 191 3791
rect 269 3589 330 3650
rect -84 2961 -23 2967
rect -84 2900 -29 2961
rect -29 2900 -23 2961
rect -84 2894 -23 2900
rect 2110 3730 2171 3791
rect 2349 3589 2410 3650
rect 2404 3305 2456 3357
rect 3595 3305 3647 3357
rect 1924 3184 1976 3236
rect 1667 3104 1719 3156
rect 269 2900 330 2961
rect 3754 3294 3806 3346
rect 3754 3184 3806 3236
rect 2404 3105 2456 3157
rect 3964 3044 4016 3096
rect 854 2750 906 2756
rect 854 2710 860 2750
rect 860 2710 900 2750
rect 900 2710 906 2750
rect 854 2704 906 2710
rect 1924 2704 1976 2756
rect 2024 2762 2088 2768
rect 2024 2698 2030 2762
rect 2030 2698 2088 2762
rect 2024 2692 2088 2698
rect 1454 2571 1506 2580
rect 1454 2537 1463 2571
rect 1463 2537 1497 2571
rect 1497 2537 1506 2571
rect 1454 2528 1506 2537
rect 2504 2528 2556 2580
rect 2634 2574 2686 2580
rect 2634 2534 2640 2574
rect 2640 2534 2680 2574
rect 2680 2534 2686 2574
rect 2634 2528 2686 2534
rect 1084 2394 1136 2446
rect 1824 2394 1876 2446
rect 2504 2404 2556 2456
rect 3964 2404 4016 2456
rect -1427 1972 -1372 2027
rect -90 1430 -30 1490
rect -688 1341 -629 1400
rect 330 1341 389 1400
rect 1830 1430 1890 1490
rect 1174 1204 1246 1276
rect 3464 1204 3536 1276
rect 6974 3294 7026 3346
rect 5374 3044 5426 3096
rect 4954 1204 5026 1276
rect 5648 1204 5720 1276
rect 6414 1204 6486 1276
rect 7248 1204 7320 1276
<< metal2 >>
rect 130 3791 191 3797
rect 191 3730 2110 3791
rect 2171 3730 2177 3791
rect 130 3724 191 3730
rect 2349 3650 2410 3656
rect 263 3589 269 3650
rect 330 3589 2349 3650
rect 2349 3583 2410 3589
rect 2404 3357 2456 3363
rect 3589 3347 3595 3357
rect 2456 3315 3595 3347
rect 3589 3305 3595 3315
rect 3647 3305 3653 3357
rect 6974 3346 7026 3352
rect 2404 3299 2456 3305
rect 3748 3294 3754 3346
rect 3806 3339 3812 3346
rect 3806 3301 6974 3339
rect 3806 3294 3812 3301
rect 6974 3288 7026 3294
rect 3754 3236 3806 3242
rect 1918 3184 1924 3236
rect 1976 3229 1982 3236
rect 1976 3191 3754 3229
rect 1976 3184 1982 3191
rect 3754 3178 3806 3184
rect 1667 3156 1719 3162
rect 2398 3147 2404 3157
rect 1719 3114 2404 3147
rect 2398 3105 2404 3114
rect 2456 3105 2462 3157
rect 1667 3098 1719 3104
rect 3964 3096 4016 3102
rect 5368 3086 5374 3096
rect 4016 3054 5374 3086
rect 5368 3044 5374 3054
rect 5426 3044 5432 3096
rect 3964 3038 4016 3044
rect -84 2967 -23 2973
rect -23 2900 269 2961
rect 330 2900 336 2961
rect -84 2888 -23 2894
rect 2024 2768 2088 2774
rect 1924 2756 1976 2762
rect 848 2704 854 2756
rect 906 2749 912 2756
rect 906 2711 1924 2749
rect 906 2704 912 2711
rect 1976 2711 2024 2749
rect 1924 2698 1976 2704
rect 2024 2686 2088 2692
rect 1454 2580 1506 2586
rect 2504 2580 2556 2586
rect 1506 2538 2504 2570
rect 1454 2522 1506 2528
rect 2628 2570 2634 2580
rect 2556 2538 2634 2570
rect 2628 2528 2634 2538
rect 2686 2528 2692 2580
rect 2504 2522 2556 2528
rect 2504 2456 2556 2462
rect 1824 2446 1876 2452
rect 1078 2394 1084 2446
rect 1136 2436 1142 2446
rect 1136 2404 1824 2436
rect 1136 2394 1142 2404
rect 3958 2446 3964 2456
rect 2556 2414 3964 2446
rect 3958 2404 3964 2414
rect 4016 2404 4022 2456
rect 2504 2398 2556 2404
rect 1824 2388 1876 2394
rect -4768 2328 -4711 2334
rect -6034 2271 -6028 2328
rect -5971 2271 -4768 2328
rect -4768 2265 -4711 2271
rect -1427 2027 -1372 2033
rect -5153 1972 -5147 2027
rect -5092 1972 -1427 2027
rect -1427 1966 -1372 1972
rect -96 1430 -90 1490
rect -30 1430 1830 1490
rect 1890 1430 1896 1490
rect -694 1341 -688 1400
rect -629 1341 330 1400
rect 389 1341 395 1400
rect 3464 1276 3536 1282
rect 6414 1276 6486 1282
rect 1168 1204 1174 1276
rect 1246 1204 3464 1276
rect 4948 1204 4954 1276
rect 5026 1204 5648 1276
rect 5720 1204 5726 1276
rect 6486 1204 7248 1276
rect 7320 1204 7326 1276
rect 3464 1198 3536 1204
rect 6414 1198 6486 1204
use CNRATR_NCH_2C8F0  CNRATR_NCH_2C8F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1709900514
transform 0 1 1124 -1 0 1236
box -184 -124 1336 1592
use CNRATR_NCH_2C8F0  CNRATR_NCH_2C8F0_1
timestamp 1709900514
transform 0 1 -376 -1 0 1236
box -184 -124 1336 1592
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -2416 -1 0 1236
box -184 -124 1336 2168
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform -1 0 6008 0 -1 3488
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_1
timestamp 1695852000
transform -1 0 7608 0 -1 2288
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_2
timestamp 1695852000
transform -1 0 6008 0 -1 4088
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_3
timestamp 1695852000
transform -1 0 7608 0 -1 3488
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_4
timestamp 1695852000
transform -1 0 7608 0 -1 4088
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_5
timestamp 1695852000
transform -1 0 7608 0 -1 4688
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_6
timestamp 1695852000
transform -1 0 6008 0 -1 2888
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_7
timestamp 1695852000
transform -1 0 7608 0 -1 2888
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_8
timestamp 1695852000
transform -1 0 6008 0 -1 2288
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_9
timestamp 1695852000
transform -1 0 6008 0 -1 4688
box -184 -124 1528 728
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 4254 -1 0 1428
box -184 -124 1528 1592
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_1
timestamp 1695852000
transform 0 1 2774 -1 0 1428
box -184 -124 1528 1592
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_2
timestamp 1695852000
transform 0 1 5714 -1 0 1428
box -184 -124 1528 1592
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_4
timestamp 1695852000
transform 0 1 -5476 -1 0 1428
box -184 -124 1528 1592
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_5
timestamp 1695852000
transform 0 1 -4016 -1 0 1428
box -184 -124 1528 1592
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_6
timestamp 1695852000
transform 0 1 -6936 -1 0 1428
box -184 -124 1528 1592
use CNRATR_NCH_8C2F0  CNRATR_NCH_8C2F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -956 -1 0 3392
box -184 -124 1912 728
use CNRATR_NCH_8C2F0  CNRATR_NCH_8C2F0_1
timestamp 1695852000
transform 0 1 -356 -1 0 3392
box -184 -124 1912 728
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 1174 -1 0 3338
box -184 -124 1528 728
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_1
timestamp 1695852000
transform 0 1 1764 -1 0 3338
box -184 -124 1528 728
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_2
timestamp 1695852000
transform 0 1 2354 -1 0 3338
box -184 -124 1528 728
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_3
timestamp 1695852000
transform 0 1 584 -1 0 3338
box -184 -124 1528 728
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -6436 -1 0 3188
box -184 -124 1528 1016
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_1
timestamp 1695852000
transform 0 1 -5556 -1 0 3188
box -184 -124 1528 1016
use CNRATR_PCH_4C12F0  CNRATR_PCH_4C12F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -4676 -1 0 3188
box -184 -124 1528 2168
use CNRATR_PCH_8C8F0  CNRATR_PCH_8C8F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -1516 -1 0 5692
box -184 -124 1912 1592
use CNRATR_PCH_8C8F0  CNRATR_PCH_8C8F0_1
timestamp 1695852000
transform 0 1 1404 -1 0 5692
box -184 -124 1912 1592
use CNRATR_PCH_8C8F0  CNRATR_PCH_8C8F0_2
timestamp 1695852000
transform 0 1 2884 -1 0 5692
box -184 -124 1912 1592
use CNRATR_PCH_8C8F0  CNRATR_PCH_8C8F0_3
timestamp 1695852000
transform 0 1 -56 -1 0 5692
box -184 -124 1912 1592
