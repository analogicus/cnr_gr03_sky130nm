magic
tech sky130B
magscale 1 2
timestamp 1713520352
<< locali >>
rect 11919 32558 20593 32559
rect 11854 32141 20593 32558
rect 11854 31592 12054 32141
rect 15219 30823 15474 30831
rect 12213 30405 19675 30823
rect 19257 23579 19675 30405
rect 20175 24405 20593 32141
rect 20175 23987 25621 24405
rect 19257 23161 25000 23579
rect 24582 22274 25000 23161
rect 25203 21871 25621 23987
rect 24582 8901 25000 10282
rect 25208 9856 28715 10274
rect 24582 8483 27893 8901
rect 422 4960 622 5346
rect 27475 4960 27893 8483
rect 422 4760 18469 4960
rect 18669 4760 27942 4960
rect 28297 4600 28715 9856
rect 27332 4400 29546 4600
rect 29346 3726 29546 4400
rect 30346 3726 30546 4160
rect 29346 3526 30558 3726
<< viali >>
rect 13326 21670 13390 21734
<< metal1 >>
rect 13320 21734 13396 21746
rect 13534 21734 13598 21740
rect 13320 21670 13326 21734
rect 13390 21670 13534 21734
rect 13320 21658 13396 21670
rect 13534 21664 13598 21670
rect 23918 19612 23924 19676
rect 23988 19612 23994 19676
rect 22900 19248 22964 19356
rect 23924 19292 23988 19612
rect 23452 19184 23458 19248
rect 23522 19184 23528 19248
rect 22900 19178 22964 19184
rect 23458 18936 23522 19184
rect 23452 18872 23458 18936
rect 23522 18872 23528 18936
<< via1 >>
rect 13534 21670 13598 21734
rect 23924 19612 23988 19676
rect 22900 19184 22964 19248
rect 23458 19184 23522 19248
rect 23458 18872 23522 18936
<< metal2 >>
rect 13733 29620 13742 29684
rect 13806 29620 13815 29684
rect 13534 21734 13598 21743
rect 13528 21670 13534 21734
rect 13598 21670 13604 21734
rect 13534 21661 13598 21670
rect 13332 21588 13396 21597
rect 13396 21524 13506 21588
rect 13332 21515 13396 21524
rect 23924 19676 23988 19682
rect 23523 19612 23532 19676
rect 23596 19612 23924 19676
rect 23924 19606 23988 19612
rect 23458 19248 23522 19254
rect 22894 19184 22900 19248
rect 22964 19184 23458 19248
rect 23458 19178 23522 19184
rect 23458 18936 23522 18942
rect 23522 18872 23702 18936
rect 23766 18872 23775 18936
rect 23458 18866 23522 18872
rect 15996 18306 16060 18310
rect 15991 18250 16000 18306
rect 16056 18250 16065 18306
rect 15996 18206 16060 18250
rect 15995 18109 16060 18206
rect 7314 8704 7378 8713
rect 7314 8631 7378 8640
rect 22705 6352 22714 6356
rect 22268 6300 22714 6352
rect 22770 6352 22779 6356
rect 22770 6300 22792 6352
rect 22268 6288 22792 6300
rect 6899 5096 6908 5152
rect 6964 5096 6973 5152
<< via2 >>
rect 13742 29620 13806 29684
rect 13534 21670 13598 21734
rect 13332 21524 13396 21588
rect 23532 19612 23596 19676
rect 23702 18872 23766 18936
rect 16000 18250 16056 18306
rect 7314 8640 7378 8704
rect 22714 6300 22770 6356
rect 6908 5096 6964 5152
<< metal3 >>
rect 16512 29816 16576 29822
rect 13736 29750 13742 29814
rect 13806 29750 13812 29814
rect 13742 29689 13806 29750
rect 13737 29684 13811 29689
rect 13737 29620 13742 29684
rect 13806 29620 13811 29684
rect 13737 29615 13811 29620
rect 16512 22242 16576 29752
rect 16506 22178 16512 22242
rect 16576 22178 16582 22242
rect 22896 22178 22902 22242
rect 22966 22178 22972 22242
rect 13529 21734 13603 21739
rect 13529 21670 13534 21734
rect 13598 21670 13603 21734
rect 13529 21665 13603 21670
rect 13327 21588 13401 21593
rect 13327 21524 13332 21588
rect 13396 21524 13401 21588
rect 13327 21519 13401 21524
rect 13332 11342 13396 21519
rect 6898 11278 6904 11342
rect 6968 11278 6974 11342
rect 13326 11278 13332 11342
rect 13396 11278 13402 11342
rect 6904 5157 6968 11278
rect 7314 11148 7378 11154
rect 13534 11148 13598 21665
rect 22902 19676 22966 22178
rect 23527 19676 23601 19681
rect 22902 19612 23532 19676
rect 23596 19612 23601 19676
rect 22902 19610 22966 19612
rect 23527 19607 23601 19612
rect 23697 18936 23771 18941
rect 23697 18872 23702 18936
rect 23766 18872 23988 18936
rect 23697 18867 23771 18872
rect 15995 18310 16061 18311
rect 15920 18306 16061 18310
rect 15920 18250 16000 18306
rect 16056 18250 16061 18306
rect 15920 18246 16061 18250
rect 15995 18245 16061 18246
rect 13528 11084 13534 11148
rect 13598 11084 13604 11148
rect 7314 8709 7378 11084
rect 7309 8704 7383 8709
rect 7309 8640 7314 8704
rect 7378 8640 7383 8704
rect 7309 8635 7383 8640
rect 23924 8172 23988 18872
rect 22704 8108 22710 8172
rect 22774 8108 22780 8172
rect 23918 8108 23924 8172
rect 23988 8108 23994 8172
rect 22710 6361 22774 8108
rect 22709 6356 22775 6361
rect 22709 6300 22714 6356
rect 22770 6300 22775 6356
rect 22709 6295 22775 6300
rect 6903 5152 6969 5157
rect 6903 5096 6908 5152
rect 6964 5096 6969 5152
rect 6903 5091 6969 5096
<< via3 >>
rect 13742 29750 13806 29814
rect 16512 29752 16576 29816
rect 16512 22178 16576 22242
rect 22902 22178 22966 22242
rect 6904 11278 6968 11342
rect 13332 11278 13396 11342
rect 7314 11084 7378 11148
rect 13534 11084 13598 11148
rect 22710 8108 22774 8172
rect 23924 8108 23988 8172
<< metal4 >>
rect 16511 29816 16577 29817
rect 13741 29814 13807 29815
rect 16511 29814 16512 29816
rect 13741 29750 13742 29814
rect 13806 29752 16512 29814
rect 16576 29814 16577 29816
rect 16576 29752 16602 29814
rect 13806 29750 16602 29752
rect 13741 29749 13807 29750
rect 16511 22242 16577 22243
rect 22901 22242 22967 22243
rect 16511 22178 16512 22242
rect 16576 22178 22902 22242
rect 22966 22178 22967 22242
rect 16511 22177 16577 22178
rect 22901 22177 22967 22178
rect 6903 11342 6969 11343
rect 13331 11342 13397 11343
rect 6903 11278 6904 11342
rect 6968 11278 13332 11342
rect 13396 11278 13397 11342
rect 6903 11277 6969 11278
rect 13331 11277 13397 11278
rect 7313 11148 7379 11149
rect 13533 11148 13599 11149
rect 7288 11084 7314 11148
rect 7378 11084 13534 11148
rect 13598 11084 13599 11148
rect 7313 11083 7379 11084
rect 13533 11083 13599 11084
rect 22709 8172 22775 8173
rect 23923 8172 23989 8173
rect 22709 8108 22710 8172
rect 22774 8108 23924 8172
rect 23988 8108 23989 8172
rect 22709 8107 22775 8108
rect 23923 8107 23989 8108
use BIAS  BIAS_0 ~/aicex/ip/cnr_gr03_sky130nm/design/CNR_GR03_SKY130NM
timestamp 1712936012
transform 0 -1 24208 1 0 15392
box -6520 -1418 7312 4136
use MILESTONE1  MILESTONE1_0
timestamp 1712303455
transform 1 0 -12348 0 1 4600
box 12340 -4600 39920 6836
use MILESTONE2  MILESTONE2_0
timestamp 1712303529
transform 0 1 11862 -1 0 30098
box -5400 -11400 18492 7028
<< labels >>
flabel locali 29346 3526 29546 4600 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel locali 422 4760 622 5346 0 FreeSans 800 0 0 0 VSS
port 2 nsew
flabel metal2 15995 18044 16060 18206 0 FreeSans 800 0 0 0 VOUT
port 3 nsew
<< end >>
