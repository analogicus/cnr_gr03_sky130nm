magic
tech sky130B
magscale 1 2
timestamp 1713190937
<< locali >>
rect 422 4960 622 5346
rect 422 4760 18469 4960
rect 18669 4760 30184 4960
rect 27332 4400 29546 4600
rect 29346 3726 29546 4400
rect 30346 3726 30546 4160
rect 29346 3526 30558 3726
<< viali >>
rect 13326 21670 13390 21734
<< metal1 >>
rect 15316 30660 15380 30666
rect 15316 30242 15380 30596
rect 15310 30178 15316 30242
rect 15380 30178 15386 30242
rect 13320 21734 13396 21746
rect 13534 21734 13598 21740
rect 13320 21670 13326 21734
rect 13390 21670 13534 21734
rect 13320 21658 13396 21670
rect 13534 21664 13598 21670
rect 22902 19356 22966 19362
rect 22902 19286 22966 19292
rect 23924 19356 23988 19362
rect 23924 19286 23988 19292
<< via1 >>
rect 15316 30596 15380 30660
rect 15316 30178 15380 30242
rect 13534 21670 13598 21734
rect 22902 19292 22966 19356
rect 23924 19292 23988 19356
<< metal2 >>
rect 15310 30596 15316 30660
rect 15380 30596 21284 30660
rect 15316 30242 15380 30248
rect 15311 30182 15316 30238
rect 15380 30182 15385 30238
rect 15316 30172 15380 30178
rect 13733 29620 13742 29684
rect 13806 29620 13815 29684
rect 15044 27202 15080 27276
rect 15023 27142 15032 27202
rect 15092 27142 15101 27202
rect 13534 21734 13598 21743
rect 13528 21670 13534 21734
rect 13598 21670 13604 21734
rect 13534 21661 13598 21670
rect 13332 21588 13396 21597
rect 13396 21524 13506 21588
rect 13332 21515 13396 21524
rect 22902 19530 22966 19539
rect 22902 19356 22966 19466
rect 22896 19292 22902 19356
rect 22966 19292 22972 19356
rect 23918 19292 23924 19356
rect 23988 19292 23994 19356
rect 23924 19174 23988 19292
rect 23924 19101 23988 19110
rect 15996 18306 16060 18310
rect 15991 18250 16000 18306
rect 16056 18250 16065 18306
rect 15996 18206 16060 18250
rect 15995 18088 16060 18206
rect 16248 18088 16312 18097
rect 15995 18045 16248 18088
rect 15996 18024 16248 18045
rect 16248 18015 16312 18024
rect 7314 8704 7378 8713
rect 7314 8631 7378 8640
rect 27036 8474 27356 8510
rect 22705 6352 22714 6356
rect 22268 6300 22714 6352
rect 22770 6352 22779 6356
rect 22770 6300 22792 6352
rect 22268 6288 22792 6300
rect 6899 5096 6908 5152
rect 6964 5096 6973 5152
<< via2 >>
rect 15320 30182 15376 30238
rect 13742 29620 13806 29684
rect 15032 27142 15092 27202
rect 13534 21670 13598 21734
rect 13332 21524 13396 21588
rect 22902 19466 22966 19530
rect 23924 19110 23988 19174
rect 16000 18250 16056 18306
rect 16248 18024 16312 18088
rect 7314 8640 7378 8704
rect 22714 6300 22770 6356
rect 6908 5096 6964 5152
<< metal3 >>
rect 15315 30238 15381 30243
rect 15315 30182 15320 30238
rect 15376 30182 15381 30238
rect 15315 30177 15381 30182
rect 15316 30012 15380 30177
rect 15310 29948 15316 30012
rect 15380 29948 15386 30012
rect 16242 29948 16248 30012
rect 16312 29948 16318 30012
rect 13736 29750 13742 29814
rect 13806 29750 13812 29814
rect 13742 29689 13806 29750
rect 13737 29684 13811 29689
rect 13737 29620 13742 29684
rect 13806 29620 13811 29684
rect 13737 29615 13811 29620
rect 15027 27202 15097 27207
rect 15027 27142 15032 27202
rect 15092 27142 15097 27202
rect 15027 27137 15097 27142
rect 15032 26996 15092 27137
rect 15024 26932 15030 26996
rect 15094 26932 15100 26996
rect 13529 21734 13603 21739
rect 13529 21670 13534 21734
rect 13598 21670 13603 21734
rect 13529 21665 13603 21670
rect 13327 21588 13401 21593
rect 13327 21524 13332 21588
rect 13396 21524 13401 21588
rect 13327 21519 13401 21524
rect 13332 11342 13396 21519
rect 6898 11278 6904 11342
rect 6968 11278 6974 11342
rect 13326 11278 13332 11342
rect 13396 11278 13402 11342
rect 6904 5157 6968 11278
rect 7314 11148 7378 11154
rect 13534 11148 13598 21665
rect 15995 18310 16061 18311
rect 15920 18306 16061 18310
rect 15920 18250 16000 18306
rect 16056 18250 16061 18306
rect 15920 18246 16061 18250
rect 15995 18245 16061 18246
rect 16248 18093 16312 29948
rect 16512 29816 16576 29822
rect 16512 22242 16576 29752
rect 17150 26932 17156 26996
rect 17220 26932 17226 26996
rect 17158 24542 17218 26932
rect 21209 24542 21329 24910
rect 17150 24478 17156 24542
rect 17220 24478 17226 24542
rect 21209 24478 21244 24542
rect 21308 24478 21329 24542
rect 21209 24414 21329 24478
rect 16506 22178 16512 22242
rect 16576 22178 16582 22242
rect 22896 22178 22902 22242
rect 22966 22178 22972 22242
rect 22902 19535 22966 22178
rect 22897 19530 22971 19535
rect 22897 19466 22902 19530
rect 22966 19466 22971 19530
rect 22897 19461 22971 19466
rect 23919 19174 23993 19179
rect 23919 19110 23924 19174
rect 23988 19110 23993 19174
rect 23919 19105 23993 19110
rect 16243 18088 16317 18093
rect 16243 18024 16248 18088
rect 16312 18024 16317 18088
rect 16243 18019 16317 18024
rect 13528 11084 13534 11148
rect 13598 11084 13604 11148
rect 7314 8709 7378 11084
rect 7309 8704 7383 8709
rect 7309 8640 7314 8704
rect 7378 8640 7383 8704
rect 7309 8635 7383 8640
rect 23924 8172 23988 19105
rect 22704 8108 22710 8172
rect 22774 8108 22780 8172
rect 23918 8108 23924 8172
rect 23988 8108 23994 8172
rect 22710 6361 22774 8108
rect 22709 6356 22775 6361
rect 22709 6300 22714 6356
rect 22770 6300 22775 6356
rect 22709 6295 22775 6300
rect 6903 5152 6969 5157
rect 6903 5096 6908 5152
rect 6964 5096 6969 5152
rect 6903 5091 6969 5096
<< via3 >>
rect 15316 29948 15380 30012
rect 16248 29948 16312 30012
rect 13742 29750 13806 29814
rect 15030 26932 15094 26996
rect 6904 11278 6968 11342
rect 13332 11278 13396 11342
rect 16512 29752 16576 29816
rect 17156 26932 17220 26996
rect 17156 24478 17220 24542
rect 21244 24478 21308 24542
rect 16512 22178 16576 22242
rect 22902 22178 22966 22242
rect 7314 11084 7378 11148
rect 13534 11084 13598 11148
rect 22710 8108 22774 8172
rect 23924 8108 23988 8172
<< metal4 >>
rect 15315 30012 15381 30013
rect 16247 30012 16313 30013
rect 15315 29948 15316 30012
rect 15380 29948 16248 30012
rect 16312 29948 16313 30012
rect 15315 29947 15381 29948
rect 16247 29947 16313 29948
rect 16511 29816 16577 29817
rect 13741 29814 13807 29815
rect 16511 29814 16512 29816
rect 13741 29750 13742 29814
rect 13806 29752 16512 29814
rect 16576 29814 16577 29816
rect 16576 29752 16602 29814
rect 13806 29750 16602 29752
rect 13741 29749 13807 29750
rect 15029 26996 15095 26997
rect 15029 26932 15030 26996
rect 15094 26994 15095 26996
rect 17155 26996 17221 26997
rect 17155 26994 17156 26996
rect 15094 26934 17156 26994
rect 15094 26932 15095 26934
rect 15029 26931 15095 26932
rect 17155 26932 17156 26934
rect 17220 26932 17221 26996
rect 17155 26931 17221 26932
rect 17155 24542 17221 24543
rect 17155 24478 17156 24542
rect 17220 24540 17221 24542
rect 21243 24542 21309 24543
rect 21243 24540 21244 24542
rect 17220 24480 21244 24540
rect 17220 24478 17221 24480
rect 17155 24477 17221 24478
rect 21243 24478 21244 24480
rect 21308 24478 21309 24542
rect 21243 24477 21309 24478
rect 16511 22242 16577 22243
rect 22901 22242 22967 22243
rect 16511 22178 16512 22242
rect 16576 22178 22902 22242
rect 22966 22178 22967 22242
rect 16511 22177 16577 22178
rect 22901 22177 22967 22178
rect 6903 11342 6969 11343
rect 13331 11342 13397 11343
rect 6903 11278 6904 11342
rect 6968 11278 13332 11342
rect 13396 11278 13397 11342
rect 6903 11277 6969 11278
rect 13331 11277 13397 11278
rect 7313 11148 7379 11149
rect 13533 11148 13599 11149
rect 7288 11084 7314 11148
rect 7378 11084 13534 11148
rect 13598 11084 13599 11148
rect 7313 11083 7379 11084
rect 13533 11083 13599 11084
rect 22709 8172 22775 8173
rect 23923 8172 23989 8173
rect 22709 8108 22710 8172
rect 22774 8108 23924 8172
rect 23988 8108 23989 8172
rect 22709 8107 22775 8108
rect 23923 8107 23989 8108
use BIAS  BIAS_0 ~/aicex/ip/cnr_gr03_sky130nm/design/CNR_GR03_SKY130NM
timestamp 1712936012
transform 0 -1 24208 1 0 15392
box -6520 -1418 7312 4136
use M3  M3_0 ~/aicex/ip/cnr_gr03_sky130nm/design/CNR_GR03_SKY130NM
timestamp 1712935398
transform 0 -1 27457 1 0 24790
box 0 2128 10317 12461
use MILESTONE1  MILESTONE1_0
timestamp 1712303455
transform 1 0 -12348 0 1 4600
box 12340 -4600 39920 6836
use MILESTONE2  MILESTONE2_0
timestamp 1712303529
transform 0 1 11862 -1 0 30098
box -5400 -11400 18492 7028
<< labels >>
flabel metal2 27036 8474 27356 8510 0 FreeSans 800 0 0 0 VRST
port 4 nsew
flabel locali 29346 3526 29546 4600 0 FreeSans 800 0 0 0 VDD
port 1 nsew
flabel locali 422 4760 622 5346 0 FreeSans 800 0 0 0 VSS
port 2 nsew
flabel space 15995 18045 16059 18251 0 FreeSans 800 180 0 0 VOUT
port 3 nsew
<< end >>
