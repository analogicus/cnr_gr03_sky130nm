magic
tech sky130B
magscale 1 2
timestamp 1712302962
<< locali >>
rect -950 5392 -584 5464
rect 650 5392 1056 5464
rect 2290 5392 2696 5464
rect 4980 4802 5016 4804
rect -2332 4557 -2177 4643
rect 657 4557 808 4643
rect -2332 4034 -2246 4557
rect -1014 4343 -777 4376
rect -743 4343 -488 4376
rect -1014 4312 -488 4343
rect 722 4063 808 4557
rect 908 4577 1043 4663
rect 3917 4617 4068 4703
rect 908 4063 994 4577
rect 2226 4312 2752 4376
rect -878 3977 -637 4063
rect 722 4034 994 4063
rect 722 3977 983 4034
rect 2362 3977 2603 4063
rect 3982 4034 4068 4617
rect 4617 4477 4703 4694
rect 4954 4358 5016 4802
rect 6600 4798 6636 4802
rect 6237 4457 6323 4694
rect 4980 4350 5016 4358
rect 6572 4362 6636 4798
rect 6572 4350 6608 4362
rect 4980 4058 5016 4062
rect 4617 3737 4703 3954
rect 4952 3622 5016 4058
rect 6572 4058 6608 4062
rect 6237 3737 6323 3954
rect 4952 3610 4988 3622
rect 6572 3622 6636 4058
rect 6600 3610 6636 3622
rect 4980 3318 5016 3322
rect 6600 3318 6636 3322
rect 1806 3084 2936 3156
rect 1806 2948 1878 3084
rect 2864 2964 2936 3084
rect 4617 2977 4703 3214
rect 4952 3148 5016 3318
rect 4952 2882 5016 3084
rect 6237 2977 6323 3214
rect 6572 3142 6636 3318
rect 6572 3090 6582 3142
rect 6634 3090 6636 3142
rect 6572 2882 6636 3090
rect 4952 2870 4988 2882
rect 6572 2870 6608 2882
rect -3786 2788 -3384 2860
rect -2746 2784 -2324 2856
rect -4138 2508 -3828 2572
rect -1470 2508 -1352 2572
rect -1288 2508 -1168 2572
rect -4592 2377 -4437 2463
rect -4592 1814 -4506 2377
rect -3892 2156 -3828 2508
rect -3892 2092 -3632 2156
rect -3568 2092 -3328 2156
rect -3892 2088 -3828 2092
rect -1232 2088 -1168 2508
rect 2548 2452 2612 2732
rect 3588 2452 3652 2592
rect 4952 2578 4988 2582
rect 6572 2578 6608 2582
rect -523 2357 -376 2443
rect 2548 2388 3652 2452
rect -3714 1737 -3477 1823
rect -2674 1737 -2417 1823
rect -462 1814 -376 2357
rect 1770 2288 2218 2316
rect 2510 2306 2958 2316
rect 1770 2280 2222 2288
rect 1782 2252 2222 2280
rect 2510 2254 2734 2306
rect 2786 2254 2958 2306
rect 2510 2252 2958 2254
rect 3250 2252 3698 2316
rect 4617 2237 4703 2474
rect 4952 2142 5016 2578
rect 6237 2237 6323 2474
rect 4980 2130 5016 2142
rect 6572 2142 6636 2578
rect 6600 2130 6636 2142
rect 250 1966 718 1976
rect 250 1948 474 1966
rect 242 1914 474 1948
rect 526 1948 718 1966
rect 526 1914 722 1948
rect 242 1912 722 1914
rect 1878 1917 2123 2003
rect 2618 1917 2843 2003
rect 3358 1917 3603 2003
rect 358 1577 603 1663
rect -6150 1068 -5764 1140
rect -4550 1068 -4184 1140
rect 4030 1062 4402 1134
rect 5630 1064 6036 1136
rect -2936 876 -2574 948
rect 830 876 1196 948
rect -6792 788 -6488 852
rect -7532 617 -7377 703
rect -7532 94 -7446 617
rect -6552 388 -6488 788
rect -2943 617 -2792 703
rect -1717 692 -1631 783
rect -1717 628 -1552 692
rect -1488 628 -926 692
rect -763 637 -616 723
rect -1717 617 -1631 628
rect -6232 372 -5668 436
rect -4632 372 -4398 436
rect -4334 372 -4068 436
rect -2878 143 -2792 617
rect -990 372 -926 628
rect -6078 57 -5857 143
rect -5518 0 -5426 80
rect -4478 57 -4257 143
rect -2878 57 -2657 143
rect -702 123 -616 637
rect 2648 637 2803 723
rect 4031 681 4188 767
rect -392 372 -328 552
rect 1206 372 1270 552
rect 2648 123 2734 637
rect -702 37 -477 123
rect 902 37 1123 123
rect 2502 94 2734 123
rect 4102 123 4188 681
rect 7243 645 7388 731
rect 4286 426 4478 436
rect 4286 374 4314 426
rect 4366 374 4478 426
rect 4286 372 4478 374
rect 5528 372 6092 436
rect 4288 328 4366 372
rect 2502 37 2723 94
rect 4102 37 4323 123
rect 5702 37 5923 123
rect 7302 94 7388 645
rect -6070 -540 -4980 0
rect -120 -540 960 10
rect 6010 -540 7100 0
rect -7100 -543 8200 -540
rect -7100 -563 6300 -543
rect -7100 -637 4680 -563
rect 4754 -617 6300 -563
rect 6374 -617 8200 -543
rect 4754 -637 8200 -617
rect -7100 -740 8200 -637
rect -7100 -963 8200 -900
rect -7100 -974 -226 -963
rect -7100 -1026 -3126 -974
rect -3074 -1026 -2206 -974
rect -2154 -1026 -226 -974
rect -7100 -1037 -226 -1026
rect -152 -1037 1294 -963
rect 1368 -1037 8200 -963
rect -7100 -1100 8200 -1037
<< viali >>
rect 8 5112 72 5176
rect 5656 5070 5720 5134
rect 7276 5038 7340 5102
rect -1586 4914 -1534 4966
rect 1654 4934 1706 4986
rect 5368 4912 5432 4976
rect 6988 4910 7052 4974
rect 3268 4728 3332 4792
rect -777 4343 -743 4377
rect 1134 4314 1186 4366
rect -2212 3928 -2148 3992
rect 7268 4386 7340 4458
rect 5368 4170 5432 4234
rect 6988 4176 7052 4240
rect 5648 3954 5720 4026
rect 5656 3568 5720 3632
rect 7268 3646 7340 3718
rect 5368 3430 5432 3494
rect 6988 3434 7052 3498
rect 74 3014 126 3066
rect 834 3014 886 3066
rect 2154 2954 2206 3006
rect 3274 2954 3326 3006
rect 4952 3084 5016 3148
rect 6582 3090 6634 3142
rect 7264 2906 7336 2978
rect 1590 2668 1654 2732
rect -3086 2514 -3034 2566
rect -1352 2508 -1288 2572
rect 80 2520 120 2560
rect 846 2513 899 2566
rect 2334 2534 2386 2586
rect -3632 2092 -3568 2156
rect 3074 2674 3126 2726
rect 3810 2668 3874 2732
rect 5368 2698 5432 2762
rect 6988 2690 7052 2754
rect -3132 1708 -3068 1772
rect 2734 2254 2786 2306
rect 5646 2474 5718 2546
rect 5656 2102 5720 2166
rect 7268 2166 7340 2238
rect 474 1914 526 1966
rect 1288 1868 1374 1954
rect 5368 1952 5432 2016
rect 6988 1958 7052 2022
rect 4974 1834 5026 1886
rect 5644 1734 5716 1806
rect 7264 1734 7336 1806
rect -232 1528 -146 1614
rect 4674 1648 4760 1734
rect 6294 1648 6380 1734
rect -5186 954 -5134 1006
rect 4990 950 5050 1010
rect 6590 950 6650 1010
rect -3586 794 -3534 846
rect 203 783 237 817
rect 1794 754 1846 806
rect 2440 800 2480 840
rect 3388 788 3452 852
rect -1552 628 -1488 692
rect -4398 372 -4334 436
rect 2892 370 2944 422
rect 4314 374 4366 426
rect 4680 -637 4754 -563
rect 6300 -617 6374 -543
rect -3126 -1026 -3074 -974
rect -2206 -1026 -2154 -974
rect -226 -1037 -152 -963
rect 1294 -1037 1368 -963
<< metal1 >>
rect 2 5182 78 5188
rect 2 5176 14 5182
rect 2 5112 8 5176
rect 2 5106 14 5112
rect 78 5106 84 5182
rect 2148 5176 2212 5182
rect 2 5100 78 5106
rect 1648 4992 1712 4998
rect -1592 4972 -1528 4978
rect -1592 4902 -1528 4908
rect -352 4972 -288 4978
rect 1302 4928 1308 4992
rect 1372 4928 1378 4992
rect -352 4512 -288 4908
rect -358 4448 -352 4512
rect -288 4448 -282 4512
rect 62 4448 68 4512
rect 132 4448 138 4512
rect -783 4377 -737 4389
rect -783 4343 -777 4377
rect -743 4343 -737 4377
rect -783 4331 -737 4343
rect -2224 3992 -2136 3998
rect -2224 3928 -2212 3992
rect -2148 3928 -2136 3992
rect -2224 3922 -2136 3928
rect -3092 2572 -3028 2578
rect -3092 2502 -3028 2508
rect -3644 2156 -3556 2162
rect -3644 2092 -3632 2156
rect -3568 2092 -3556 2156
rect -3644 2086 -3556 2092
rect -3632 1672 -3568 2086
rect -3144 1772 -3056 1778
rect -3144 1708 -3132 1772
rect -3068 1708 -3056 1772
rect -3144 1702 -3056 1708
rect -5198 1608 -5192 1672
rect -5128 1608 -5122 1672
rect -5192 1006 -5128 1608
rect -3632 1602 -3568 1608
rect -5192 954 -5186 1006
rect -5134 954 -5128 1006
rect -5192 942 -5128 954
rect -3592 852 -3528 858
rect -3592 782 -3528 788
rect -4410 436 -4322 442
rect -4410 372 -4398 436
rect -4334 372 -4322 436
rect -4410 366 -4322 372
rect -4398 322 -4334 366
rect -4398 252 -4334 258
rect -3132 -974 -3068 1702
rect -2398 1628 -2392 1692
rect -2328 1628 -2322 1692
rect -2392 852 -2328 1628
rect -2398 788 -2392 852
rect -2328 788 -2322 852
rect -2212 -968 -2148 3922
rect -782 3792 -738 4331
rect -786 3786 -734 3792
rect -786 3728 -734 3734
rect -386 3786 -334 3792
rect -386 3728 -334 3734
rect -1364 2572 -1276 2578
rect -1558 2508 -1552 2572
rect -1488 2508 -1482 2572
rect -1364 2508 -1352 2572
rect -1288 2508 -1276 2572
rect -382 2566 -338 3728
rect 68 3072 132 4448
rect 1128 4366 1192 4378
rect 1128 4314 1134 4366
rect 1186 4314 1192 4366
rect 828 3840 892 3846
rect 62 3066 138 3072
rect 62 3014 74 3066
rect 126 3014 138 3066
rect 62 3008 138 3014
rect 828 3066 892 3776
rect 828 3014 834 3066
rect 886 3014 892 3066
rect 828 3002 892 3014
rect 74 2566 126 2572
rect -392 2514 -386 2566
rect -334 2514 -328 2566
rect -1552 1572 -1488 2508
rect -1364 2502 -1276 2508
rect -1352 1692 -1288 2502
rect -1352 1622 -1288 1628
rect -1558 1508 -1552 1572
rect -1488 1508 -1482 1572
rect -1552 698 -1488 1508
rect -382 1072 -338 2514
rect 74 2508 126 2514
rect 840 2566 905 2578
rect 840 2513 846 2566
rect 899 2513 905 2566
rect 468 1966 532 1978
rect 468 1914 474 1966
rect 526 1914 532 1966
rect 468 1692 532 1914
rect 840 1840 905 2513
rect 1128 2232 1192 4314
rect 1308 3840 1372 4928
rect 1648 4922 1712 4928
rect 1308 3770 1372 3776
rect 2148 3006 2212 5112
rect 5650 5140 5726 5146
rect 5650 5134 5662 5140
rect 5650 5070 5656 5134
rect 5650 5064 5662 5070
rect 5726 5064 5732 5140
rect 5976 5134 6040 5140
rect 7270 5108 7346 5114
rect 5650 5058 5726 5064
rect 5362 4982 5438 4988
rect 5362 4976 5374 4982
rect 5362 4912 5368 4976
rect 5362 4906 5374 4912
rect 5438 4906 5444 4982
rect 5758 4912 5764 4976
rect 5828 4912 5834 4976
rect 5362 4900 5438 4906
rect 3256 4792 3344 4798
rect 3256 4728 3268 4792
rect 3332 4728 3344 4792
rect 3256 4722 3344 4728
rect 3268 3012 3332 4722
rect 5362 4290 5368 4354
rect 5432 4290 5438 4354
rect 5368 4246 5432 4290
rect 5764 4246 5828 4912
rect 5976 4464 6040 5070
rect 6248 5102 6312 5108
rect 5976 4458 6050 4464
rect 5976 4386 5978 4458
rect 5976 4380 6050 4386
rect 5362 4234 5438 4246
rect 5362 4170 5368 4234
rect 5432 4170 5438 4234
rect 5362 4158 5438 4170
rect 5764 4240 5832 4246
rect 5764 4176 5768 4240
rect 5764 4170 5832 4176
rect 5642 4032 5726 4038
rect 5642 4026 5654 4032
rect 5642 3954 5648 4026
rect 5642 3948 5654 3954
rect 5726 3948 5732 4032
rect 5642 3942 5726 3948
rect 5650 3638 5726 3644
rect 5650 3632 5662 3638
rect 5650 3568 5656 3632
rect 5650 3562 5662 3568
rect 5726 3562 5732 3638
rect 5650 3556 5726 3562
rect 5362 3500 5438 3506
rect 5362 3494 5374 3500
rect 5362 3430 5368 3494
rect 5362 3424 5374 3430
rect 5438 3424 5444 3500
rect 5764 3494 5828 4170
rect 5362 3418 5438 3424
rect 4946 3154 5022 3160
rect 4946 3148 4958 3154
rect 4946 3084 4952 3148
rect 4946 3078 4958 3084
rect 5022 3078 5028 3154
rect 4946 3072 5022 3078
rect 2148 2954 2154 3006
rect 2206 2954 2212 3006
rect 2148 2942 2212 2954
rect 3262 3006 3338 3012
rect 3262 2954 3274 3006
rect 3326 2954 3338 3006
rect 5764 2998 5828 3430
rect 5976 3638 6040 4380
rect 6248 4032 6312 5038
rect 7264 5032 7270 5108
rect 7334 5102 7346 5108
rect 7340 5038 7346 5102
rect 7334 5032 7346 5038
rect 7270 5026 7346 5032
rect 6982 4980 7058 4986
rect 6432 4910 6438 4974
rect 6502 4910 6508 4974
rect 6438 4354 6502 4910
rect 6976 4904 6982 4980
rect 7046 4974 7058 4980
rect 7052 4910 7058 4974
rect 7046 4904 7058 4910
rect 6982 4898 7058 4904
rect 7262 4464 7346 4470
rect 7256 4380 7262 4464
rect 7334 4458 7346 4464
rect 7340 4386 7346 4458
rect 7334 4380 7346 4386
rect 7262 4374 7346 4380
rect 6242 4026 6314 4032
rect 6242 3948 6314 3954
rect 6248 3724 6312 3948
rect 6248 3718 6324 3724
rect 6248 3646 6252 3718
rect 6248 3640 6324 3646
rect 5976 3632 6044 3638
rect 5976 3568 5980 3632
rect 5976 3562 6044 3568
rect 3262 2948 3338 2954
rect 4790 2934 4796 2998
rect 4860 2934 4866 2998
rect 5758 2934 5764 2998
rect 5828 2934 5834 2998
rect 5976 2984 6040 3562
rect 5976 2978 6048 2984
rect 1584 2738 1660 2744
rect 1584 2732 1596 2738
rect 1584 2668 1590 2732
rect 1584 2662 1596 2668
rect 1660 2662 1666 2738
rect 3068 2732 3132 2738
rect 3068 2662 3132 2668
rect 3804 2732 3880 2744
rect 4796 2734 4860 2934
rect 5362 2796 5368 2860
rect 5432 2796 5438 2860
rect 5368 2768 5432 2796
rect 3804 2668 3810 2732
rect 3874 2668 3880 2732
rect 4302 2668 4308 2732
rect 4372 2668 4378 2732
rect 5356 2762 5444 2768
rect 5356 2698 5368 2762
rect 5432 2698 5444 2762
rect 5356 2692 5444 2698
rect 5764 2754 5828 2934
rect 1584 2656 1660 2662
rect 3804 2656 3880 2668
rect 2328 2586 2392 2598
rect 2328 2534 2334 2586
rect 2386 2534 2392 2586
rect 2328 2472 2392 2534
rect 2328 2402 2392 2408
rect 3810 2472 3874 2656
rect 3810 2402 3874 2408
rect 840 1834 913 1840
rect 840 1769 848 1834
rect 840 1763 913 1769
rect 1127 1834 1192 2232
rect 2728 2306 2792 2318
rect 2728 2254 2734 2306
rect 2786 2254 2792 2306
rect 1276 1954 1386 1960
rect 1276 1868 1288 1954
rect 1374 1868 1386 1954
rect 1276 1862 1386 1868
rect 1127 1763 1192 1769
rect 462 1628 468 1692
rect 532 1628 538 1692
rect -244 1614 -134 1620
rect -244 1528 -232 1614
rect -146 1528 -134 1614
rect -244 1522 -134 1528
rect -386 1066 -334 1072
rect -386 1008 -334 1014
rect -1564 692 -1476 698
rect -1564 628 -1552 692
rect -1488 628 -1476 692
rect -1564 622 -1476 628
rect -232 -963 -146 1522
rect 840 1072 905 1763
rect 194 1066 246 1072
rect 194 1008 246 1014
rect 834 1008 840 1072
rect 904 1008 910 1072
rect 198 829 242 1008
rect 197 817 243 829
rect 197 783 203 817
rect 237 783 243 817
rect 197 771 243 783
rect 1288 -957 1374 1862
rect 2728 1692 2792 2254
rect 2728 1622 2792 1628
rect 1782 1008 1788 1072
rect 1852 1008 1858 1072
rect 1788 806 1852 1008
rect 3382 858 3458 864
rect 1788 754 1794 806
rect 1846 754 1852 806
rect 2434 846 2486 852
rect 2434 788 2486 794
rect 3376 782 3382 858
rect 3434 852 3458 858
rect 3452 788 3458 852
rect 3434 782 3458 788
rect 3382 776 3458 782
rect 1788 742 1852 754
rect 2886 422 2950 434
rect 2886 370 2892 422
rect 2944 370 2950 422
rect 2886 322 2950 370
rect 4308 426 4372 2668
rect 4796 2664 4860 2670
rect 5640 2552 5724 2558
rect 5640 2546 5652 2552
rect 4402 2472 4466 2478
rect 5640 2474 5646 2546
rect 5640 2468 5652 2474
rect 5724 2468 5730 2552
rect 5640 2462 5724 2468
rect 4402 2362 4466 2408
rect 4402 2292 4466 2298
rect 5650 2172 5726 2178
rect 5650 2166 5662 2172
rect 5650 2102 5656 2166
rect 5650 2096 5662 2102
rect 5726 2096 5732 2172
rect 5650 2090 5726 2096
rect 5362 2022 5438 2028
rect 5362 2016 5374 2022
rect 5362 1952 5368 2016
rect 5362 1946 5374 1952
rect 5438 1946 5444 2022
rect 5764 2016 5828 2690
rect 5976 2900 6048 2906
rect 5976 2166 6040 2900
rect 6248 2552 6312 3640
rect 6438 3498 6502 4290
rect 6982 4246 7058 4252
rect 6976 4170 6982 4246
rect 7046 4240 7058 4246
rect 7052 4176 7058 4240
rect 7046 4170 7058 4176
rect 6982 4164 7058 4170
rect 7262 3724 7346 3730
rect 7256 3640 7262 3724
rect 7334 3718 7346 3724
rect 7340 3646 7346 3718
rect 7334 3640 7346 3646
rect 7262 3634 7346 3640
rect 6982 3504 7058 3510
rect 6438 2866 6502 3434
rect 6976 3428 6982 3504
rect 7046 3498 7058 3504
rect 7052 3434 7058 3498
rect 7046 3428 7058 3434
rect 6982 3422 7058 3428
rect 6576 3148 6640 3154
rect 6576 3078 6640 3084
rect 7258 2984 7342 2990
rect 7252 2900 7258 2984
rect 7330 2978 7342 2984
rect 7336 2906 7342 2978
rect 7330 2900 7342 2906
rect 7258 2894 7342 2900
rect 6438 2860 6506 2866
rect 6438 2796 6442 2860
rect 6438 2790 6506 2796
rect 6242 2546 6314 2552
rect 6242 2468 6314 2474
rect 6248 2244 6312 2468
rect 6438 2362 6502 2790
rect 6982 2760 7058 2766
rect 6976 2684 6982 2760
rect 7046 2754 7058 2760
rect 7052 2690 7058 2754
rect 7046 2684 7058 2690
rect 6982 2678 7058 2684
rect 6432 2298 6438 2362
rect 6502 2298 6508 2362
rect 6248 2238 6324 2244
rect 6248 2166 6252 2238
rect 6248 2160 6324 2166
rect 6248 2102 6312 2160
rect 5976 2094 6040 2102
rect 5764 1946 5828 1952
rect 6438 2028 6502 2298
rect 7262 2244 7346 2250
rect 7256 2160 7262 2244
rect 7334 2238 7346 2244
rect 7340 2166 7346 2238
rect 7334 2160 7346 2166
rect 7262 2154 7346 2160
rect 6982 2028 7058 2034
rect 6438 2022 6506 2028
rect 6438 1958 6442 2022
rect 6438 1952 6506 1958
rect 6976 1952 6982 2028
rect 7046 2022 7058 2028
rect 7052 1958 7058 2022
rect 7046 1952 7058 1958
rect 6438 1948 6502 1952
rect 6982 1946 7058 1952
rect 5362 1940 5438 1946
rect 4968 1886 5032 1898
rect 4968 1834 4974 1886
rect 5026 1834 5032 1886
rect 4662 1734 4772 1740
rect 4662 1648 4674 1734
rect 4760 1648 4772 1734
rect 4662 1642 4772 1648
rect 4308 374 4314 426
rect 4366 374 4372 426
rect 4308 362 4372 374
rect 2886 252 2950 258
rect 4674 -563 4760 1642
rect 4968 1572 5032 1834
rect 5632 1806 5728 1812
rect 5632 1734 5644 1806
rect 5716 1734 5728 1806
rect 7252 1806 7348 1812
rect 5632 1728 5728 1734
rect 6282 1734 6392 1740
rect 4962 1508 4968 1572
rect 5032 1508 5038 1572
rect 5644 1276 5716 1728
rect 6282 1648 6294 1734
rect 6380 1648 6392 1734
rect 7252 1734 7264 1806
rect 7336 1734 7348 1806
rect 7252 1728 7348 1734
rect 6282 1642 6392 1648
rect 4978 1204 4984 1276
rect 5056 1204 5062 1276
rect 4984 1010 5056 1204
rect 5644 1198 5716 1204
rect 4984 950 4990 1010
rect 5050 950 5056 1010
rect 4984 938 5056 950
rect 4674 -637 4680 -563
rect 4754 -637 4760 -563
rect 6294 -543 6380 1642
rect 7264 1276 7336 1728
rect 6578 1204 6584 1276
rect 6656 1204 6662 1276
rect 6584 1010 6656 1204
rect 7264 1198 7336 1204
rect 6584 950 6590 1010
rect 6650 950 6656 1010
rect 6584 938 6656 950
rect 6294 -617 6300 -543
rect 6374 -617 6380 -543
rect 6294 -629 6380 -617
rect 4674 -649 4760 -637
rect -3132 -1026 -3126 -974
rect -3074 -1026 -3068 -974
rect -3132 -1038 -3068 -1026
rect -2218 -974 -2142 -968
rect -2218 -1026 -2206 -974
rect -2154 -1026 -2142 -974
rect -2218 -1032 -2142 -1026
rect -232 -1037 -226 -963
rect -152 -1037 -146 -963
rect -232 -1049 -146 -1037
rect 1282 -963 1380 -957
rect 1282 -1037 1294 -963
rect 1368 -1037 1380 -963
rect 1282 -1043 1380 -1037
<< via1 >>
rect 14 5176 78 5182
rect 14 5112 72 5176
rect 72 5112 78 5176
rect 14 5106 78 5112
rect 2148 5112 2212 5176
rect -1592 4966 -1528 4972
rect -1592 4914 -1586 4966
rect -1586 4914 -1534 4966
rect -1534 4914 -1528 4966
rect -1592 4908 -1528 4914
rect -352 4908 -288 4972
rect 1308 4928 1372 4992
rect 1648 4986 1712 4992
rect 1648 4934 1654 4986
rect 1654 4934 1706 4986
rect 1706 4934 1712 4986
rect 1648 4928 1712 4934
rect -352 4448 -288 4512
rect 68 4448 132 4512
rect -3092 2566 -3028 2572
rect -3092 2514 -3086 2566
rect -3086 2514 -3034 2566
rect -3034 2514 -3028 2566
rect -3092 2508 -3028 2514
rect -5192 1608 -5128 1672
rect -3632 1608 -3568 1672
rect -3592 846 -3528 852
rect -3592 794 -3586 846
rect -3586 794 -3534 846
rect -3534 794 -3528 846
rect -3592 788 -3528 794
rect -4398 258 -4334 322
rect -2392 1628 -2328 1692
rect -2392 788 -2328 852
rect -786 3734 -734 3786
rect -386 3734 -334 3786
rect -1552 2508 -1488 2572
rect 828 3776 892 3840
rect -386 2514 -334 2566
rect 74 2560 126 2566
rect 74 2520 80 2560
rect 80 2520 120 2560
rect 120 2520 126 2560
rect 74 2514 126 2520
rect -1352 1628 -1288 1692
rect -1552 1508 -1488 1572
rect 1308 3776 1372 3840
rect 5662 5134 5726 5140
rect 5662 5070 5720 5134
rect 5720 5070 5726 5134
rect 5662 5064 5726 5070
rect 5976 5070 6040 5134
rect 5374 4976 5438 4982
rect 5374 4912 5432 4976
rect 5432 4912 5438 4976
rect 5374 4906 5438 4912
rect 5764 4912 5828 4976
rect 5368 4290 5432 4354
rect 6248 5038 6312 5102
rect 5978 4386 6050 4458
rect 5768 4176 5832 4240
rect 5654 4026 5726 4032
rect 5654 3954 5720 4026
rect 5720 3954 5726 4026
rect 5654 3948 5726 3954
rect 5662 3632 5726 3638
rect 5662 3568 5720 3632
rect 5720 3568 5726 3632
rect 5662 3562 5726 3568
rect 5374 3494 5438 3500
rect 5374 3430 5432 3494
rect 5432 3430 5438 3494
rect 5374 3424 5438 3430
rect 5764 3430 5828 3494
rect 4958 3148 5022 3154
rect 4958 3084 5016 3148
rect 5016 3084 5022 3148
rect 4958 3078 5022 3084
rect 7270 5102 7334 5108
rect 7270 5038 7276 5102
rect 7276 5038 7334 5102
rect 7270 5032 7334 5038
rect 6438 4910 6502 4974
rect 6982 4974 7046 4980
rect 6982 4910 6988 4974
rect 6988 4910 7046 4974
rect 6982 4904 7046 4910
rect 7262 4458 7334 4464
rect 7262 4386 7268 4458
rect 7268 4386 7334 4458
rect 7262 4380 7334 4386
rect 6438 4290 6502 4354
rect 6242 3954 6314 4026
rect 6252 3646 6324 3718
rect 5980 3568 6044 3632
rect 4796 2934 4860 2998
rect 5764 2934 5828 2998
rect 1596 2732 1660 2738
rect 1596 2668 1654 2732
rect 1654 2668 1660 2732
rect 1596 2662 1660 2668
rect 3068 2726 3132 2732
rect 3068 2674 3074 2726
rect 3074 2674 3126 2726
rect 3126 2674 3132 2726
rect 3068 2668 3132 2674
rect 5368 2796 5432 2860
rect 4308 2668 4372 2732
rect 4796 2670 4860 2734
rect 2328 2408 2392 2472
rect 3810 2408 3874 2472
rect 848 1769 913 1834
rect 1127 1769 1192 1834
rect 468 1628 532 1692
rect -386 1014 -334 1066
rect 194 1014 246 1066
rect 840 1008 904 1072
rect 2728 1628 2792 1692
rect 1788 1008 1852 1072
rect 2434 840 2486 846
rect 2434 800 2440 840
rect 2440 800 2480 840
rect 2480 800 2486 840
rect 2434 794 2486 800
rect 3382 852 3434 858
rect 3382 788 3388 852
rect 3388 788 3434 852
rect 3382 782 3434 788
rect 5764 2690 5828 2754
rect 5652 2546 5724 2552
rect 4402 2408 4466 2472
rect 5652 2474 5718 2546
rect 5718 2474 5724 2546
rect 5652 2468 5724 2474
rect 4402 2298 4466 2362
rect 5662 2166 5726 2172
rect 5662 2102 5720 2166
rect 5720 2102 5726 2166
rect 5662 2096 5726 2102
rect 5374 2016 5438 2022
rect 5374 1952 5432 2016
rect 5432 1952 5438 2016
rect 5374 1946 5438 1952
rect 5976 2906 6048 2978
rect 6982 4240 7046 4246
rect 6982 4176 6988 4240
rect 6988 4176 7046 4240
rect 6982 4170 7046 4176
rect 7262 3718 7334 3724
rect 7262 3646 7268 3718
rect 7268 3646 7334 3718
rect 7262 3640 7334 3646
rect 6438 3434 6502 3498
rect 6982 3498 7046 3504
rect 6982 3434 6988 3498
rect 6988 3434 7046 3498
rect 6982 3428 7046 3434
rect 6576 3142 6640 3148
rect 6576 3090 6582 3142
rect 6582 3090 6634 3142
rect 6634 3090 6640 3142
rect 6576 3084 6640 3090
rect 7258 2978 7330 2984
rect 7258 2906 7264 2978
rect 7264 2906 7330 2978
rect 7258 2900 7330 2906
rect 6442 2796 6506 2860
rect 6242 2474 6314 2546
rect 5976 2102 6040 2166
rect 6982 2754 7046 2760
rect 6982 2690 6988 2754
rect 6988 2690 7046 2754
rect 6982 2684 7046 2690
rect 6438 2298 6502 2362
rect 6252 2166 6324 2238
rect 5764 1952 5828 2016
rect 7262 2238 7334 2244
rect 7262 2166 7268 2238
rect 7268 2166 7334 2238
rect 7262 2160 7334 2166
rect 6442 1958 6506 2022
rect 6982 2022 7046 2028
rect 6982 1958 6988 2022
rect 6988 1958 7046 2022
rect 6982 1952 7046 1958
rect 2886 258 2950 322
rect 4968 1508 5032 1572
rect 4984 1204 5056 1276
rect 5644 1204 5716 1276
rect 6584 1204 6656 1276
rect 7264 1204 7336 1276
<< metal2 >>
rect 14 5182 78 5188
rect 78 5112 2148 5176
rect 2212 5112 2218 5176
rect 5662 5140 5726 5146
rect 14 5100 78 5106
rect 5726 5070 5976 5134
rect 6040 5070 6046 5134
rect 7270 5108 7334 5114
rect 5662 5058 5726 5064
rect 6242 5038 6248 5102
rect 6312 5038 7270 5102
rect 7270 5026 7334 5032
rect 1308 4992 1372 4998
rect -1598 4908 -1592 4972
rect -1528 4908 -352 4972
rect -288 4908 -280 4972
rect 1300 4928 1308 4992
rect 1372 4928 1648 4992
rect 1712 4928 1718 4992
rect 5374 4982 5438 4988
rect 1308 4922 1372 4928
rect 5764 4976 5828 4982
rect 6982 4980 7046 4986
rect 5438 4912 5764 4976
rect 5764 4906 5828 4912
rect 6438 4974 6502 4980
rect 6502 4910 6982 4974
rect 5374 4900 5438 4906
rect 6438 4904 6502 4910
rect 6982 4898 7046 4904
rect -352 4512 -288 4518
rect 68 4512 132 4518
rect -288 4448 68 4512
rect 7262 4464 7334 4470
rect -352 4442 -288 4448
rect 68 4442 132 4448
rect 5972 4386 5978 4458
rect 6050 4386 7262 4458
rect 7262 4374 7334 4380
rect 5368 4354 5432 4360
rect 5432 4290 6438 4354
rect 6502 4290 6508 4354
rect 5368 4284 5432 4290
rect 6982 4246 7046 4252
rect 5762 4176 5768 4240
rect 5832 4176 6982 4240
rect 6982 4164 7046 4170
rect 5654 4032 5726 4038
rect 5726 3954 6242 4026
rect 6314 3954 6320 4026
rect 5654 3942 5726 3948
rect -792 3734 -786 3786
rect -734 3782 -728 3786
rect -392 3782 -386 3786
rect -734 3738 -386 3782
rect -734 3734 -728 3738
rect -392 3734 -386 3738
rect -334 3734 -328 3786
rect 822 3776 828 3840
rect 892 3776 1308 3840
rect 1372 3776 1378 3840
rect 7262 3724 7334 3730
rect 6246 3646 6252 3718
rect 6324 3646 7262 3718
rect 5662 3638 5726 3644
rect 7262 3634 7334 3640
rect 5726 3568 5980 3632
rect 6044 3568 6050 3632
rect 5662 3556 5726 3562
rect 5374 3500 5438 3506
rect 6982 3504 7046 3510
rect 5438 3430 5764 3494
rect 5828 3430 5834 3494
rect 6432 3434 6438 3498
rect 6502 3434 6982 3498
rect 5374 3418 5438 3424
rect 6982 3422 7046 3428
rect 4958 3154 5022 3160
rect 5022 3084 6576 3148
rect 6640 3084 6646 3148
rect 4958 3072 5022 3078
rect 4796 2998 4860 3004
rect 5764 2998 5828 3004
rect 4860 2934 5764 2998
rect 7258 2984 7330 2990
rect 4796 2928 4860 2934
rect 5764 2928 5828 2934
rect 5970 2906 5976 2978
rect 6048 2906 7258 2978
rect 7258 2894 7330 2900
rect 5368 2860 5432 2866
rect 5432 2796 6442 2860
rect 6506 2796 6512 2860
rect 5368 2790 5432 2796
rect 6982 2760 7046 2766
rect 1596 2738 1660 2744
rect 4308 2732 4372 2738
rect 4790 2732 4796 2734
rect 1660 2668 3068 2732
rect 3132 2668 4308 2732
rect 4372 2670 4796 2732
rect 4860 2670 4866 2734
rect 5758 2690 5764 2754
rect 5828 2690 6982 2754
rect 6982 2678 7046 2684
rect 4372 2668 4866 2670
rect 4308 2662 4372 2668
rect 1596 2656 1660 2662
rect -1552 2572 -1488 2578
rect -3098 2508 -3092 2572
rect -3028 2508 -1552 2572
rect -386 2566 -334 2572
rect 68 2562 74 2566
rect -334 2518 74 2562
rect 68 2514 74 2518
rect 126 2514 132 2566
rect 5652 2552 5724 2558
rect -386 2508 -334 2514
rect -1552 2502 -1488 2508
rect 2322 2408 2328 2472
rect 2392 2408 3810 2472
rect 3874 2408 4402 2472
rect 4466 2408 4472 2472
rect 5724 2474 6242 2546
rect 6314 2474 6320 2546
rect 5652 2462 5724 2468
rect 6438 2362 6502 2368
rect 4396 2298 4402 2362
rect 4466 2298 6438 2362
rect 6438 2292 6502 2298
rect 7262 2244 7334 2250
rect 5662 2172 5726 2178
rect 6246 2166 6252 2238
rect 6324 2166 7262 2238
rect 5726 2102 5976 2166
rect 6040 2102 6046 2166
rect 7262 2154 7334 2160
rect 5662 2090 5726 2096
rect 6982 2028 7046 2034
rect 5374 2022 5438 2028
rect 5438 1952 5764 2016
rect 5828 1952 5834 2016
rect 6436 1958 6442 2022
rect 6506 1958 6982 2022
rect 6982 1946 7046 1952
rect 5374 1940 5438 1946
rect 842 1769 848 1834
rect 913 1769 1127 1834
rect 1192 1769 1198 1834
rect -2392 1692 -2328 1698
rect 468 1692 532 1698
rect -5192 1672 -5128 1678
rect -5128 1608 -3632 1672
rect -3568 1608 -3562 1672
rect -2328 1628 -1352 1692
rect -1288 1628 468 1692
rect 532 1628 2728 1692
rect 2792 1628 2798 1692
rect -2392 1622 -2328 1628
rect 468 1622 532 1628
rect -5192 1602 -5128 1608
rect -1552 1572 -1488 1578
rect 4968 1572 5032 1578
rect -1488 1508 4968 1572
rect -1552 1502 -1488 1508
rect 4968 1502 5032 1508
rect 4984 1276 5056 1282
rect 6584 1276 6656 1282
rect 5056 1204 5644 1276
rect 5716 1204 5722 1276
rect 6656 1204 7264 1276
rect 7336 1204 7342 1276
rect 4984 1198 5056 1204
rect 6584 1198 6656 1204
rect 840 1072 904 1078
rect 1788 1072 1852 1078
rect -392 1014 -386 1066
rect -334 1062 -328 1066
rect 188 1062 194 1066
rect -334 1018 194 1062
rect -334 1014 -328 1018
rect 188 1014 194 1018
rect 246 1014 252 1066
rect 904 1008 1788 1072
rect 840 1002 904 1008
rect 1788 1002 1852 1008
rect 3382 858 3434 864
rect -2392 852 -2328 858
rect -3598 788 -3592 852
rect -3528 788 -2392 852
rect 2428 794 2434 846
rect 2486 794 3382 846
rect -2392 782 -2328 788
rect 3382 776 3434 782
rect -4404 258 -4398 322
rect -4334 258 2886 322
rect 2950 258 2956 322
use CNRATR_NCH_2C8F0  CNRATR_NCH_2C8F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1709900514
transform 0 1 1084 -1 0 1236
box -184 -124 1336 1592
use CNRATR_NCH_2C8F0  CNRATR_NCH_2C8F0_1
timestamp 1709900514
transform 0 1 -516 -1 0 1236
box -184 -124 1336 1592
use CNRATR_NCH_2C12F0  CNRATR_NCH_2C12F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -2696 -1 0 1236
box -184 -124 1336 2168
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform -1 0 6008 0 -1 3768
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_1
timestamp 1695852000
transform -1 0 7628 0 -1 2288
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_2
timestamp 1695852000
transform -1 0 6008 0 -1 4508
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_3
timestamp 1695852000
transform -1 0 7628 0 -1 3768
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_4
timestamp 1695852000
transform -1 0 7628 0 -1 4508
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_5
timestamp 1695852000
transform -1 0 7628 0 -1 5248
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_6
timestamp 1695852000
transform -1 0 6008 0 -1 3028
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_7
timestamp 1695852000
transform -1 0 7628 0 -1 3028
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_8
timestamp 1695852000
transform -1 0 6008 0 -1 2288
box -184 -124 1528 728
use CNRATR_NCH_4C2F0  CNRATR_NCH_4C2F0_9
timestamp 1695852000
transform -1 0 6008 0 -1 5248
box -184 -124 1528 728
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 4284 -1 0 1428
box -184 -124 1528 1592
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_1
timestamp 1695852000
transform 0 1 2684 -1 0 1428
box -184 -124 1528 1592
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_2
timestamp 1695852000
transform 0 1 5884 -1 0 1428
box -184 -124 1528 1592
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_4
timestamp 1695852000
transform 0 1 -5896 -1 0 1428
box -184 -124 1528 1592
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_5
timestamp 1695852000
transform 0 1 -4296 -1 0 1428
box -184 -124 1528 1592
use CNRATR_NCH_4C8F0  CNRATR_NCH_4C8F0_6
timestamp 1695852000
transform 0 1 -7496 -1 0 1428
box -184 -124 1528 1592
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 2064 -1 0 3308
box -184 -124 1528 728
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_1
timestamp 1695852000
transform 0 1 2804 -1 0 3308
box -184 -124 1528 728
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_2
timestamp 1695852000
transform 0 1 3544 -1 0 3308
box -184 -124 1528 728
use CNRATR_PCH_4C2F0  CNRATR_PCH_4C2F0_3
timestamp 1695852000
transform 0 1 1324 -1 0 3308
box -184 -124 1528 728
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -4556 -1 0 3148
box -184 -124 1528 1016
use CNRATR_PCH_4C4F0  CNRATR_PCH_4C4F0_1
timestamp 1695852000
transform 0 1 -3516 -1 0 3148
box -184 -124 1528 1016
use CNRATR_PCH_4C12F0  CNRATR_PCH_4C12F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -2456 -1 0 3148
box -184 -124 1528 2168
use CNRATR_PCH_8C2F0  CNRATR_PCH_8C2F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -196 -1 0 3352
box -184 -124 1912 728
use CNRATR_PCH_8C2F0  CNRATR_PCH_8C2F0_1
timestamp 1695852000
transform 0 1 564 -1 0 3352
box -184 -124 1912 728
use CNRATR_PCH_8C8F0  CNRATR_PCH_8C8F0_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -2296 -1 0 5752
box -184 -124 1912 1592
use CNRATR_PCH_8C8F0  CNRATR_PCH_8C8F0_1
timestamp 1695852000
transform 0 1 944 -1 0 5752
box -184 -124 1912 1592
use CNRATR_PCH_8C8F0  CNRATR_PCH_8C8F0_2
timestamp 1695852000
transform 0 1 2564 -1 0 5752
box -184 -124 1912 1592
use CNRATR_PCH_8C8F0  CNRATR_PCH_8C8F0_3
timestamp 1695852000
transform 0 1 -696 -1 0 5752
box -184 -124 1912 1592
<< labels >>
flabel locali 1368 -1100 8200 -900 0 FreeSans 800 0 0 0 VDD
port 7 nsew
flabel locali 1368 -740 4680 -540 0 FreeSans 800 0 0 0 VSS
port 10 nsew
flabel locali -6798 788 -6488 852 0 FreeSans 800 0 0 0 IBIAS
port 11 nsew
flabel locali -392 372 -328 552 0 FreeSans 800 0 0 0 VIP
port 9 nsew
flabel locali 1206 372 1270 552 0 FreeSans 800 0 0 0 VIN
port 8 nsew
flabel metal2 4466 2298 6438 2362 0 FreeSans 800 0 0 0 VOUT
port 12 nsew
<< end >>
