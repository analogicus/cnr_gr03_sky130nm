** sch_path: /home/ocheid/aicex/ip/cnr_gr03_sky130nm/design/CNR_GR03_SKY130NM/MILESTONE1.sch
**.subckt MILESTONE1 VDD VSS I_OUT1 I_OUT2
*.iopin VDD
*.iopin VSS
*.iopin I_OUT1
*.iopin I_OUT2
V0 I_OUT1 VSS 0
x3<20> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<19> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<18> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<17> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<16> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<15> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<14> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<13> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<12> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<11> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<10> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<9> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<8> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<7> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<6> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<5> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<4> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<3> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<2> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<1> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x3<0> I_OUT1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<20> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<19> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<18> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<17> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<16> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<15> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<14> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<13> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<12> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<11> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<10> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<9> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<8> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<7> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<6> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<5> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<4> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<3> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<2> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<1> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x2<0> VR1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<20> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<19> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<18> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<17> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<16> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<15> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<14> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<13> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<12> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<11> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<10> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<9> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<8> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<7> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<6> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<5> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<4> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<3> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<2> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<1> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x5<0> VD1 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
R1 VR1 VD2 1k m=1
XQ1 VSS VSS VD1 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=1
XQ2 VSS VSS VD2 sky130_fd_pr__pnp_05v5_W3p40L3p40 m=5
x1<20> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<19> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<18> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<17> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<16> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<15> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<14> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<13> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<12> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<11> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<10> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<9> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<8> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<7> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<6> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<5> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<4> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<3> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<2> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<1> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1<0> I_OUT2 OTA_OUT VDD VDD CNRATR_PCH_8C1F2
x1 VDD VR1 OTA_OUT VD1 IBIAS VSS CM_OTA_NCH
I0 VDD IBIAS 2u
**.ends

* expanding   symbol:
*+  /home/ocheid/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_8C1F2.sym # of pins=4
** sym_path: /home/ocheid/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_8C1F2.sym
** sch_path: /home/ocheid/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_8C1F2.sch
.subckt CNRATR_PCH_8C1F2 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=0.252 W=7.68 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  CNR_GR03_SKY130NM/CM_OTA_NCH.sym # of pins=6
** sym_path: /home/ocheid/aicex/ip/cnr_gr03_sky130nm/design/CNR_GR03_SKY130NM/CM_OTA_NCH.sym
** sch_path: /home/ocheid/aicex/ip/cnr_gr03_sky130nm/design/CNR_GR03_SKY130NM/CM_OTA_NCH.sch
.subckt CM_OTA_NCH VDD VIP VOUT VIN IBIAS VSS
*.iopin VDD
*.iopin VIN
*.iopin VIP
*.iopin VSS
*.iopin IBIAS
*.iopin VOUT
x13 VBP1 VIN VS VSS CNRATR_NCH_8C8F0
x1 VBP2 VIP VS VSS CNRATR_NCH_8C8F0
x2 VS IBIAS VSS VSS CNRATR_NCH_4C8F0
x3 IBIAS IBIAS VSS VSS CNRATR_NCH_4C8F0
x5 VBP1 VBP1 VDD VDD CNRATR_PCH_8C8F0
x4 Vn1 VBP1 VDD VDD CNRATR_PCH_8C8F0
x6 VBP2 VBP2 VDD VDD CNRATR_PCH_8C8F0
x7 VOUT VBP2 VDD VDD CNRATR_PCH_8C8F0
x8 Vn1 Vn1 VSS VSS CNRATR_NCH_4C8F0
x9 VOUT Vn1 VSS VSS CNRATR_NCH_4C8F0
.ends


* expanding   symbol:
*+  /home/ocheid/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_8C8F0.sym # of pins=4
** sym_path: /home/ocheid/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_8C8F0.sym
** sch_path: /home/ocheid/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_8C8F0.sch
.subckt CNRATR_NCH_8C8F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=2.7 W=7.68 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:
*+  /home/ocheid/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_4C8F0.sym # of pins=4
** sym_path: /home/ocheid/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_4C8F0.sym
** sch_path: /home/ocheid/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_NCH_4C8F0.sch
.subckt CNRATR_NCH_4C8F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__nfet_01v8 L=2.7 W=3.84 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:
*+  /home/ocheid/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_8C8F0.sym # of pins=4
** sym_path: /home/ocheid/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_8C8F0.sym
** sch_path: /home/ocheid/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM/CNRATR_PCH_8C8F0.sch
.subckt CNRATR_PCH_8C8F0 D G S B
*.iopin D
*.iopin G
*.iopin S
*.iopin B
XM1 D G S B sky130_fd_pr__pfet_01v8 L=2.7 W=7.68 nf=2 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
