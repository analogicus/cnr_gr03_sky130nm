*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/MILESTONE1_lpe.spi
#else
.include ../../../work/xsch/MILESTONE1.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15 reltol=1e-6 abstol=1e-6 keepopinfo noopiter gminsteps=5

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS VSS 0 dc 0
VDD VDD 0 dc 1.8 
IBIAS VDD IBIAS dc 2u
*V0 OTA_OUT 0 dc 0
V0 IOUT1 VSS dc 0

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD VSS IOUT1 VREF IBIAS MILESTONE1

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
.save v(VSS) v(VDD) v(XDUT.VD1) v(XDUT.VR1) v(XDUT.VD2) v(XDUT.OTA_OUT) v(IOUT1) v(VREF) i(v.XDUT.V1)
.save i(V0)

#endifmak

*----------------------------------------------------------------
* NGSPICE controlplo
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 10n 10u 0

#ifdef Debug
tran 10p 1n 1p
*quit
#else
tran 10p 10n 1p
dc temp -40 125 2 
write
quit
#endif

.endc

.end
