*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/MILESTONE2_lpe.spi
#else
.include ../../../work/xsch/MILESTONE2.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0 dc 0
VDD  VDD_1V8 VSS dc 1.8
Vrst RST VSS PULSE(0 1.8 0.0 2NS 2NS 1MS 2MS)
Iin I_IN VSS dc 1u
Vref VREF_I VSS dc 1.2

*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT RST OUT I_IN VREF_I VDD_1V8 VSS MILESTONE2

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

#ifdef Debug
.save all
#else
*.save *v(OUT)
.save all
#endif

*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

optran 0 0 0 10n 10u 0

#ifdef Debug
tran 10p 1n 1p
*quit
#else
*tran 1u 10m
tran 10p 10n 1p
dc Iin 50u 75u 100n
write
quit
#endif

.endc

.end
