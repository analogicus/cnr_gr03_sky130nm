magic
tech sky130B
magscale 1 2
timestamp 1710172682
<< locali >>
rect -9599 9712 -9344 9784
rect -9090 9710 -8814 9782
rect -8610 9720 -8355 9792
rect -8100 9710 -7824 9782
rect -7619 9712 -7364 9784
rect -7110 9710 -6834 9782
rect -6630 9720 -6375 9792
rect -6150 9720 -5874 9792
rect -5649 9712 -5394 9784
rect -5150 9720 -4874 9792
rect -4660 9720 -4405 9792
rect -4170 9710 -3894 9782
rect -3649 9712 -3394 9784
rect -3140 9720 -2864 9792
rect -2660 9710 -2405 9782
rect -2140 9720 -1864 9792
rect -1620 9710 -1344 9782
rect -1140 9720 -864 9792
rect -660 9710 -384 9782
rect -160 9720 116 9792
rect 4101 9732 4356 9804
rect 4610 9740 4886 9812
rect 5090 9740 5345 9812
rect 5590 9730 5866 9802
rect 6081 9732 6336 9804
rect 6580 9740 6856 9812
rect 7070 9740 7325 9812
rect 7560 9740 7836 9812
rect 8051 9732 8306 9804
rect 8550 9740 8826 9812
rect 9040 9740 9295 9812
rect 9520 9730 9796 9802
rect 10051 9732 10306 9804
rect 10540 9730 10816 9802
rect 11040 9730 11295 9802
rect 11580 9730 11856 9802
rect 12060 9730 12336 9802
rect 12560 9730 12836 9802
rect 13040 9730 13316 9802
rect 13540 9730 13816 9802
rect -9638 8632 -9332 8689
rect -9120 8640 -8804 8696
rect -8640 8630 -8334 8687
rect -8140 8640 -7824 8696
rect -7658 8632 -7352 8689
rect -7140 8640 -6824 8696
rect -6660 8630 -6354 8687
rect -6160 8640 -5844 8696
rect -5688 8632 -5382 8689
rect -5170 8640 -4854 8696
rect -4690 8630 -4384 8687
rect -4190 8640 -3874 8696
rect -3688 8632 -3382 8689
rect -3170 8640 -2854 8696
rect -2690 8630 -2384 8687
rect -2160 8640 -1844 8696
rect -1660 8640 -1344 8696
rect -1170 8640 -854 8696
rect -680 8640 -364 8696
rect -190 8640 126 8696
rect 4062 8652 4368 8709
rect 4562 8652 4878 8708
rect 5060 8650 5366 8707
rect 5570 8660 5886 8716
rect 6042 8652 6348 8709
rect 6570 8660 6886 8716
rect 7040 8650 7346 8707
rect 7540 8660 7856 8716
rect 8012 8652 8318 8709
rect 8530 8660 8846 8716
rect 9010 8650 9316 8707
rect 9510 8660 9826 8716
rect 10012 8652 10318 8709
rect 10530 8660 10846 8716
rect 11010 8650 11316 8707
rect 11540 8660 11856 8716
rect 12040 8660 12356 8716
rect 12530 8660 12846 8716
rect 13030 8660 13346 8716
rect 13510 8660 13826 8716
rect -9589 7322 -9334 7394
rect -9080 7330 -8804 7402
rect -8600 7330 -8345 7402
rect -8100 7320 -7824 7392
rect -7609 7322 -7354 7394
rect -7110 7330 -6834 7402
rect -6620 7330 -6365 7402
rect -6130 7330 -5854 7402
rect -5639 7322 -5384 7394
rect -5140 7330 -4864 7402
rect -4650 7330 -4395 7402
rect -4170 7320 -3894 7392
rect -3639 7322 -3384 7394
rect -3150 7320 -2874 7392
rect -2650 7320 -2395 7392
rect -2110 7320 -1834 7392
rect -1630 7320 -1354 7392
rect -1130 7320 -854 7392
rect -650 7320 -374 7392
rect -150 7320 126 7392
rect -9628 6242 -9322 6299
rect -9128 6242 -8812 6298
rect -8630 6240 -8324 6297
rect -8120 6250 -7804 6306
rect -7648 6242 -7342 6299
rect -7120 6250 -6804 6306
rect -6650 6240 -6344 6297
rect -6150 6250 -5834 6306
rect -5678 6242 -5372 6299
rect -5160 6250 -4844 6306
rect -4680 6240 -4374 6297
rect -4180 6250 -3864 6306
rect -3678 6242 -3372 6299
rect -3160 6250 -2844 6306
rect -2680 6240 -2374 6297
rect -2150 6250 -1834 6306
rect -1650 6250 -1334 6306
rect -1160 6250 -844 6306
rect -660 6250 -344 6306
rect -180 6250 136 6306
rect -10200 310 178 510
rect -10200 0 180 200
use CM_OTA_NCH  CM_OTA_NCH_0
timestamp 1710170680
transform 1 0 7078 0 1 1050
box -7100 -1050 8200 5876
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -4536 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_1
timestamp 1695852000
transform 0 1 -5026 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_2
timestamp 1695852000
transform 0 1 -5516 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_3
timestamp 1695852000
transform 0 1 -6016 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_4
timestamp 1695852000
transform 0 1 -8486 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_5
timestamp 1695852000
transform 0 1 -8976 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_6
timestamp 1695852000
transform 0 1 -9456 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_7
timestamp 1695852000
transform 0 1 -9956 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_8
timestamp 1695852000
transform 0 1 -7986 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_9
timestamp 1695852000
transform 0 1 -7486 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_10
timestamp 1695852000
transform 0 1 -6996 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_11
timestamp 1695852000
transform 0 1 -6496 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_12
timestamp 1695852000
transform 0 1 -2506 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_13
timestamp 1695852000
transform 0 1 -526 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_14
timestamp 1695852000
transform 0 1 -3026 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_15
timestamp 1695852000
transform 0 1 -2006 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_16
timestamp 1695852000
transform 0 1 -1516 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_17
timestamp 1695852000
transform 0 1 -3506 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_18
timestamp 1695852000
transform 0 1 -4006 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_19
timestamp 1695852000
transform 0 1 -1016 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_20
timestamp 1695852000
transform 0 1 -16 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_21
timestamp 1695852000
transform 0 1 -9466 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_22
timestamp 1695852000
transform 0 1 -9966 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_23
timestamp 1695852000
transform 0 1 -6986 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_24
timestamp 1695852000
transform 0 1 -7476 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_25
timestamp 1695852000
transform 0 1 -8476 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_26
timestamp 1695852000
transform 0 1 -7976 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_27
timestamp 1695852000
transform 0 1 -8966 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_28
timestamp 1695852000
transform 0 1 -6506 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_29
timestamp 1695852000
transform 0 1 -4526 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_30
timestamp 1695852000
transform 0 1 -5506 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_31
timestamp 1695852000
transform 0 1 -5016 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_32
timestamp 1695852000
transform 0 1 -6006 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_33
timestamp 1695852000
transform 0 1 -3516 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_34
timestamp 1695852000
transform 0 1 -4016 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_35
timestamp 1695852000
transform 0 1 -1506 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_36
timestamp 1695852000
transform 0 1 -2496 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_37
timestamp 1695852000
transform 0 1 -1996 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_38
timestamp 1695852000
transform 0 1 -3016 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_39
timestamp 1695852000
transform 0 1 -536 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_40
timestamp 1695852000
transform 0 1 -1026 -1 0 10072
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_41
timestamp 1695852000
transform 0 1 -6 -1 0 7682
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_42
timestamp 1695852000
transform 0 1 13684 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_43
timestamp 1695852000
transform 0 1 13164 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_44
timestamp 1695852000
transform 0 1 12674 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_45
timestamp 1695852000
transform 0 1 12184 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_46
timestamp 1695852000
transform 0 1 11694 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_47
timestamp 1695852000
transform 0 1 11194 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_48
timestamp 1695852000
transform 0 1 10674 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_49
timestamp 1695852000
transform 0 1 10184 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_50
timestamp 1695852000
transform 0 1 9684 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_51
timestamp 1695852000
transform 0 1 8674 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_52
timestamp 1695852000
transform 0 1 9164 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_53
timestamp 1695852000
transform 0 1 8184 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_54
timestamp 1695852000
transform 0 1 7684 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_55
timestamp 1695852000
transform 0 1 6704 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_56
timestamp 1695852000
transform 0 1 7194 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_57
timestamp 1695852000
transform 0 1 6214 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_58
timestamp 1695852000
transform 0 1 5714 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_59
timestamp 1695852000
transform 0 1 4724 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_60
timestamp 1695852000
transform 0 1 5214 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_61
timestamp 1695852000
transform 0 1 3734 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_62
timestamp 1695852000
transform 0 1 4234 -1 0 10092
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_63
timestamp 1695852000
transform 0 1 3534 -1 0 7602
box -184 -124 1912 613
use sky130_fd_pr__rf_pnp_05v5_W0p68L0p68  sky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1704988097
transform 1 0 -14940 0 1 2670
box 0 0 796 796
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1704988097
transform 1 0 -12110 0 1 2220
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1704988097
transform 1 0 -13880 0 1 2320
box 0 0 1340 1340
<< end >>
