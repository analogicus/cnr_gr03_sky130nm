magic
tech sky130B
magscale 1 2
timestamp 1710522302
<< locali >>
rect -6360 4794 -6304 4802
rect -7089 4722 -6824 4794
rect -6579 4730 -6304 4794
rect -6579 4722 -6344 4730
rect -6100 4720 -5824 4792
rect -5600 4730 -5324 4802
rect -5089 4722 -4314 4794
rect -4069 4722 -3814 4794
rect -3560 4730 -3284 4802
rect -3080 4730 -2825 4802
rect -2580 4720 -2328 4792
rect -2109 4722 -1354 4794
rect -7492 3977 -7317 4063
rect -7492 3364 -7406 3977
rect -7403 3907 -7317 3977
rect -2103 3887 -1951 4053
rect -7130 3650 -6813 3706
rect -6610 3650 -6293 3706
rect -6120 3653 -5804 3706
rect -6099 3650 -5804 3653
rect -5630 3650 -5314 3706
rect -5128 3642 -4262 3682
rect -4090 3650 -3774 3707
rect -3590 3650 -3274 3707
rect -3100 3650 -2784 3707
rect -2610 3650 -2498 3707
rect -2441 3650 -2328 3707
rect -2037 3453 -1951 3887
rect -5000 3260 -4400 3440
rect -2037 3297 -1427 3453
rect 7819 3381 8021 3383
rect 7819 3341 7820 3381
rect 7860 3341 8021 3381
rect 7819 3340 8021 3341
rect -1513 3277 -1427 3297
rect -307 2616 -248 2702
rect -2370 2350 -2094 2422
rect -1870 2350 -1594 2422
rect -1390 2350 -1153 2422
rect -890 2350 -614 2422
rect 5850 1768 5882 1870
rect -2772 1527 -2627 1743
rect 5830 1704 6440 1768
rect -5056 824 -4984 1061
rect -4720 510 -4520 960
rect -4411 824 -4339 1061
rect -2772 1000 -2686 1527
rect -373 1497 -221 1633
rect -2390 1280 -2074 1336
rect -1900 1327 -1584 1336
rect -1900 1293 -1785 1327
rect -1751 1293 -1584 1327
rect -1900 1280 -1584 1293
rect -1400 1280 -1084 1336
rect -921 1280 -604 1336
rect -307 1000 -221 1497
rect 6376 1424 6440 1704
rect 6838 510 6934 1134
rect 15919 1004 15991 1241
rect 16052 510 16151 1105
rect -10700 450 17780 510
rect -10700 432 6610 450
rect -10700 367 -7732 432
rect -7667 430 6610 432
rect -7667 367 -5070 430
rect -10700 330 -5070 367
rect -4970 414 6610 430
rect -4970 345 -2314 414
rect -2245 350 6610 414
rect 6710 350 17780 450
rect -2245 345 17780 350
rect -4970 330 17780 345
rect -10700 310 17780 330
rect -10700 127 18220 200
rect -10700 53 -7486 127
rect -7412 53 18220 127
rect -10700 0 18220 53
rect -5256 -492 -5076 -380
rect -4964 -492 -4864 -380
rect -2456 -461 -2336 -380
rect -2224 -461 -2084 -380
rect -2456 -492 -2084 -461
rect 6364 -492 6604 -380
rect 6716 -492 6956 -380
rect 7360 -997 7636 -942
rect 7360 -1107 7405 -997
rect 7515 -1107 7636 -997
rect 7360 -1162 7636 -1107
<< viali >>
rect 7155 5310 7205 5360
rect -7230 4259 -7190 4299
rect -6720 4259 -6680 4299
rect -6240 4259 -6200 4299
rect -5750 4259 -5710 4299
rect -5230 4259 -5190 4299
rect -4192 4250 -4156 4314
rect -3710 4262 -3670 4302
rect -3220 4262 -3180 4302
rect -2730 4262 -2690 4302
rect -2250 4262 -2210 4302
rect 6581 3981 6619 4019
rect -2498 3650 -2441 3707
rect -1243 3657 -1198 3702
rect -7492 3258 -7406 3344
rect 3599 3330 3640 3390
rect 7820 3341 7860 3381
rect 6885 3024 6919 3058
rect -2520 1892 -2480 1932
rect -2020 1892 -1980 1932
rect -1530 1892 -1490 1932
rect -1040 1892 -1000 1932
rect -520 1892 -480 1932
rect -1785 1293 -1751 1327
rect 7016 1422 7080 1486
rect 8518 1422 8582 1486
rect -7732 367 -7667 432
rect -5070 330 -4970 430
rect -2314 345 -2245 414
rect 6610 350 6710 450
rect -7486 53 -7412 127
rect -7756 -457 -7644 -380
rect -5076 -492 -4964 -380
rect -2336 -461 -2224 -380
rect 6604 -492 6716 -380
rect -6837 -1077 -6803 -1043
rect -5947 -1067 -5893 -1013
rect -3937 -1057 -3903 -1023
rect -3092 -1162 -2944 -942
rect -1588 -1120 -1452 -984
rect 5782 -1162 5904 -942
rect 7405 -1107 7515 -997
rect 14774 -1086 14826 -1034
<< metal1 >>
rect 7143 5360 7217 5366
rect 7143 5310 7155 5360
rect 7205 5310 7217 5360
rect 7143 5304 7217 5310
rect 6574 4726 6626 4732
rect 7155 4726 7205 5304
rect 7148 4674 7154 4726
rect 7206 4674 7212 4726
rect 6574 4668 6626 4674
rect -4198 4320 -4150 4326
rect -7236 4305 -7184 4311
rect -7236 4247 -7184 4253
rect -6726 4305 -6674 4311
rect -6726 4247 -6674 4253
rect -6246 4305 -6194 4311
rect -6246 4247 -6194 4253
rect -5756 4305 -5704 4311
rect -5236 4305 -5184 4311
rect -5492 4253 -5486 4305
rect -5434 4253 -5428 4305
rect -5756 4247 -5704 4253
rect -7504 3344 -7394 3350
rect -7504 3258 -7492 3344
rect -7406 3258 -7394 3344
rect -7504 3252 -7394 3258
rect -7738 432 -7661 444
rect -7738 367 -7732 432
rect -7667 367 -7661 432
rect -7738 -374 -7661 367
rect -7492 127 -7406 3252
rect -6852 3041 -6846 3093
rect -6794 3041 -6788 3093
rect -6834 2478 -6806 3041
rect -6852 2472 -6788 2478
rect -6852 2402 -6788 2408
rect -7492 53 -7486 127
rect -7412 53 -7406 127
rect -7492 41 -7406 53
rect -7768 -380 -7632 -374
rect -7768 -457 -7756 -380
rect -7644 -457 -7632 -380
rect -7768 -463 -7632 -457
rect -6834 -1031 -6806 2402
rect -5474 1886 -5446 4253
rect -5236 4247 -5184 4253
rect -4206 4244 -4200 4320
rect -4148 4244 -4142 4320
rect -3716 4308 -3664 4314
rect -3972 4256 -3966 4308
rect -3914 4256 -3908 4308
rect -4198 4238 -4150 4244
rect -3954 3099 -3926 4256
rect -3716 4250 -3664 4256
rect -3226 4308 -3174 4314
rect -2256 4308 -2204 4314
rect -2742 4256 -2736 4308
rect -2684 4256 -2678 4308
rect -3226 4250 -3174 4256
rect -2256 4250 -2204 4256
rect 6575 4019 6625 4668
rect 10526 4234 10532 4286
rect 10584 4234 10590 4286
rect 6575 3981 6581 4019
rect 6619 3981 6625 4019
rect 6575 3969 6625 3981
rect 10539 3916 10577 4234
rect 10532 3910 10584 3916
rect 10532 3852 10584 3858
rect -2510 3707 -2429 3713
rect -2510 3650 -2498 3707
rect -2441 3650 -2429 3707
rect -2510 3644 -2429 3650
rect -1589 3702 -1186 3708
rect -1589 3657 -1243 3702
rect -1198 3657 -1186 3702
rect -1589 3651 -1186 3657
rect -2497 3579 -2440 3644
rect -1589 3579 -1532 3651
rect -1805 3522 -1799 3574
rect -1738 3522 -1732 3574
rect -2497 3516 -2440 3522
rect -3966 3093 -3914 3099
rect -3966 3035 -3914 3041
rect -1791 3060 -1745 3522
rect -1589 3516 -1532 3522
rect 3593 3396 3646 3402
rect 3588 3324 3594 3396
rect 3646 3324 3652 3396
rect 7814 3387 7866 3393
rect 6869 3335 6875 3387
rect 6927 3335 6933 3387
rect 3593 3318 3646 3324
rect 6880 3070 6923 3335
rect 7814 3329 7866 3335
rect -1791 3054 -1726 3060
rect -1791 2994 -1786 3054
rect 6879 3058 6925 3070
rect 6879 3024 6885 3058
rect 6919 3024 6925 3058
rect 6879 3012 6925 3024
rect -1791 2988 -1726 2994
rect -3006 1938 -2954 1944
rect -2026 1938 -1974 1944
rect -2532 1886 -2526 1938
rect -2474 1886 -2468 1938
rect -5491 1880 -5429 1886
rect -3006 1880 -2954 1886
rect -2026 1880 -1974 1886
rect -5059 1818 -5053 1880
rect -4991 1818 -4985 1880
rect -5491 1812 -5429 1818
rect -5474 1806 -5446 1812
rect -5053 1169 -4991 1818
rect -5076 430 -4964 442
rect -5076 330 -5070 430
rect -4970 330 -4964 430
rect -5953 113 -5887 119
rect -5953 -1007 -5887 47
rect -5076 -374 -4964 330
rect -3970 113 -3904 1513
rect -3976 47 -3970 113
rect -3904 47 -3898 113
rect -2997 -128 -2963 1880
rect -1791 1333 -1745 2988
rect -1536 1938 -1484 1944
rect -1536 1880 -1484 1886
rect -1046 1938 -994 1944
rect -1046 1880 -994 1886
rect -526 1938 -474 1944
rect -526 1880 -474 1886
rect 7004 1486 7092 1492
rect 7004 1480 7016 1486
rect 7080 1480 7092 1486
rect 7004 1416 7010 1480
rect 7086 1416 7092 1480
rect 8506 1486 8594 1492
rect 8506 1480 8518 1486
rect 8582 1480 8594 1486
rect 8506 1416 8512 1480
rect 8588 1416 8594 1480
rect 7010 1410 7086 1416
rect 8512 1410 8588 1416
rect -1797 1327 -1739 1333
rect -1797 1293 -1785 1327
rect -1751 1293 -1739 1327
rect -1797 1287 -1739 1293
rect 15470 787 15536 1693
rect 6604 450 6716 462
rect -2320 414 -2239 426
rect -2320 345 -2314 414
rect -2245 345 -2239 414
rect -3006 -134 -2954 -128
rect -3952 -186 -3946 -134
rect -3894 -186 -3888 -134
rect -5088 -380 -4952 -374
rect -5088 -492 -5076 -380
rect -4964 -492 -4952 -380
rect -5088 -498 -4952 -492
rect -5959 -1013 -5881 -1007
rect -6843 -1043 -6797 -1031
rect -6843 -1077 -6837 -1043
rect -6803 -1077 -6797 -1043
rect -5959 -1067 -5947 -1013
rect -5893 -1067 -5881 -1013
rect -3937 -1017 -3903 -186
rect -3006 -192 -2954 -186
rect -2320 -374 -2239 345
rect 6604 350 6610 450
rect 6710 350 6716 450
rect 6604 -374 6716 350
rect -2348 -380 -2212 -374
rect -2348 -461 -2336 -380
rect -2224 -461 -2212 -380
rect -2348 -467 -2212 -461
rect 6592 -380 6728 -374
rect 6592 -492 6604 -380
rect 6716 -492 6728 -380
rect 6592 -498 6728 -492
rect -3098 -936 -2938 -930
rect 5776 -936 5910 -930
rect -3098 -942 -3086 -936
rect -3949 -1023 -3891 -1017
rect -3949 -1057 -3937 -1023
rect -3903 -1057 -3891 -1023
rect -3949 -1063 -3891 -1057
rect -5959 -1073 -5881 -1067
rect -6843 -1089 -6797 -1077
rect -3098 -1162 -3092 -942
rect -3098 -1168 -3086 -1162
rect -2938 -1168 -2932 -936
rect 5776 -942 5788 -936
rect -1594 -978 -1446 -972
rect -1594 -1132 -1446 -1126
rect 5776 -1162 5782 -942
rect 5776 -1168 5788 -1162
rect 5910 -1168 5916 -936
rect 7399 -991 7521 -985
rect 14768 -1028 14832 -1022
rect 15471 -1028 15535 787
rect 15465 -1092 15471 -1028
rect 15535 -1092 15541 -1028
rect 14768 -1098 14832 -1092
rect 7399 -1119 7521 -1113
rect -3098 -1174 -2938 -1168
rect 5776 -1174 5910 -1168
<< via1 >>
rect 6574 4674 6626 4726
rect 7154 4674 7206 4726
rect -7236 4299 -7184 4305
rect -7236 4259 -7230 4299
rect -7230 4259 -7190 4299
rect -7190 4259 -7184 4299
rect -7236 4253 -7184 4259
rect -6726 4299 -6674 4305
rect -6726 4259 -6720 4299
rect -6720 4259 -6680 4299
rect -6680 4259 -6674 4299
rect -6726 4253 -6674 4259
rect -6246 4299 -6194 4305
rect -6246 4259 -6240 4299
rect -6240 4259 -6200 4299
rect -6200 4259 -6194 4299
rect -6246 4253 -6194 4259
rect -5756 4299 -5704 4305
rect -5756 4259 -5750 4299
rect -5750 4259 -5710 4299
rect -5710 4259 -5704 4299
rect -5756 4253 -5704 4259
rect -5486 4253 -5434 4305
rect -5236 4299 -5184 4305
rect -5236 4259 -5230 4299
rect -5230 4259 -5190 4299
rect -5190 4259 -5184 4299
rect -5236 4253 -5184 4259
rect -6846 3041 -6794 3093
rect -6852 2408 -6788 2472
rect -4200 4314 -4148 4320
rect -4200 4250 -4192 4314
rect -4192 4250 -4156 4314
rect -4156 4250 -4148 4314
rect -4200 4244 -4148 4250
rect -3966 4256 -3914 4308
rect -3716 4302 -3664 4308
rect -3716 4262 -3710 4302
rect -3710 4262 -3670 4302
rect -3670 4262 -3664 4302
rect -3716 4256 -3664 4262
rect -3226 4302 -3174 4308
rect -3226 4262 -3220 4302
rect -3220 4262 -3180 4302
rect -3180 4262 -3174 4302
rect -3226 4256 -3174 4262
rect -2736 4302 -2684 4308
rect -2736 4262 -2730 4302
rect -2730 4262 -2690 4302
rect -2690 4262 -2684 4302
rect -2736 4256 -2684 4262
rect -2256 4302 -2204 4308
rect -2256 4262 -2250 4302
rect -2250 4262 -2210 4302
rect -2210 4262 -2204 4302
rect -2256 4256 -2204 4262
rect 10532 4234 10584 4286
rect 10532 3858 10584 3910
rect -2497 3522 -2440 3579
rect -1799 3522 -1738 3574
rect -1589 3522 -1532 3579
rect -3966 3041 -3914 3093
rect 3594 3390 3646 3396
rect 3594 3330 3599 3390
rect 3599 3330 3640 3390
rect 3640 3330 3646 3390
rect 3594 3324 3646 3330
rect 6875 3335 6927 3387
rect 7814 3381 7866 3387
rect 7814 3341 7820 3381
rect 7820 3341 7860 3381
rect 7860 3341 7866 3381
rect 7814 3335 7866 3341
rect -1786 2994 -1726 3054
rect -3006 1886 -2954 1938
rect -2526 1932 -2474 1938
rect -2526 1892 -2520 1932
rect -2520 1892 -2480 1932
rect -2480 1892 -2474 1932
rect -2526 1886 -2474 1892
rect -2026 1932 -1974 1938
rect -2026 1892 -2020 1932
rect -2020 1892 -1980 1932
rect -1980 1892 -1974 1932
rect -2026 1886 -1974 1892
rect -5491 1818 -5429 1880
rect -5053 1818 -4991 1880
rect -5953 47 -5887 113
rect -3970 47 -3904 113
rect -1536 1932 -1484 1938
rect -1536 1892 -1530 1932
rect -1530 1892 -1490 1932
rect -1490 1892 -1484 1932
rect -1536 1886 -1484 1892
rect -1046 1932 -994 1938
rect -1046 1892 -1040 1932
rect -1040 1892 -1000 1932
rect -1000 1892 -994 1932
rect -1046 1886 -994 1892
rect -526 1932 -474 1938
rect -526 1892 -520 1932
rect -520 1892 -480 1932
rect -480 1892 -474 1932
rect -526 1886 -474 1892
rect 7010 1422 7016 1480
rect 7016 1422 7080 1480
rect 7080 1422 7086 1480
rect 7010 1416 7086 1422
rect 8512 1422 8518 1480
rect 8518 1422 8582 1480
rect 8582 1422 8588 1480
rect 8512 1416 8588 1422
rect -3946 -186 -3894 -134
rect -3006 -186 -2954 -134
rect -3086 -942 -2938 -936
rect -3086 -1162 -2944 -942
rect -2944 -1162 -2938 -942
rect -3086 -1168 -2938 -1162
rect 5788 -942 5910 -936
rect -1594 -984 -1446 -978
rect -1594 -1120 -1588 -984
rect -1588 -1120 -1452 -984
rect -1452 -1120 -1446 -984
rect -1594 -1126 -1446 -1120
rect 5788 -1162 5904 -942
rect 5904 -1162 5910 -942
rect 5788 -1168 5910 -1162
rect 7399 -997 7521 -991
rect 7399 -1107 7405 -997
rect 7405 -1107 7515 -997
rect 7515 -1107 7521 -997
rect 14768 -1034 14832 -1028
rect 14768 -1086 14774 -1034
rect 14774 -1086 14826 -1034
rect 14826 -1086 14832 -1034
rect 14768 -1092 14832 -1086
rect 15471 -1092 15535 -1028
rect 7399 -1113 7521 -1107
<< metal2 >>
rect 7154 4726 7206 4732
rect 6568 4674 6574 4726
rect 6626 4725 6632 4726
rect 6626 4675 7154 4725
rect 6626 4674 6632 4675
rect 7154 4668 7206 4674
rect -4200 4320 -4148 4326
rect -5486 4305 -5434 4311
rect -7242 4253 -7236 4305
rect -7184 4297 -7178 4305
rect -6732 4297 -6726 4305
rect -7184 4261 -6726 4297
rect -7184 4253 -7178 4261
rect -6732 4253 -6726 4261
rect -6674 4297 -6668 4305
rect -6252 4297 -6246 4305
rect -6674 4261 -6246 4297
rect -6674 4253 -6668 4261
rect -6252 4253 -6246 4261
rect -6194 4297 -6188 4305
rect -5762 4297 -5756 4305
rect -6194 4261 -5756 4297
rect -6194 4253 -6188 4261
rect -5762 4253 -5756 4261
rect -5704 4297 -5698 4305
rect -5704 4261 -5486 4297
rect -5704 4253 -5698 4261
rect -5242 4297 -5236 4305
rect -5434 4261 -5236 4297
rect -5242 4253 -5236 4261
rect -5184 4253 -5178 4305
rect -5486 4247 -5434 4253
rect -3966 4308 -3914 4314
rect -2736 4308 -2684 4314
rect -4148 4264 -3966 4300
rect -3722 4300 -3716 4308
rect -3914 4264 -3716 4300
rect -3722 4256 -3716 4264
rect -3664 4300 -3658 4308
rect -3232 4300 -3226 4308
rect -3664 4264 -3226 4300
rect -3664 4256 -3658 4264
rect -3232 4256 -3226 4264
rect -3174 4300 -3168 4308
rect -3174 4264 -2736 4300
rect -3174 4256 -3168 4264
rect -2262 4300 -2256 4308
rect -2684 4264 -2256 4300
rect -2262 4256 -2256 4264
rect -2204 4256 -2198 4308
rect 10532 4286 10584 4292
rect -3966 4250 -3914 4256
rect -2736 4250 -2684 4256
rect -4200 4238 -4148 4244
rect 10532 4228 10584 4234
rect 10528 3914 10588 3923
rect 10526 3858 10528 3910
rect 10588 3858 10590 3910
rect 10528 3845 10588 3854
rect -1799 3579 -1738 3580
rect -2503 3522 -2497 3579
rect -2440 3574 -1589 3579
rect -2440 3522 -1799 3574
rect -1738 3522 -1589 3574
rect -1532 3522 -1526 3579
rect -1799 3516 -1738 3522
rect 3594 3396 3646 3402
rect 6875 3387 6927 3393
rect 3646 3339 6875 3382
rect 7808 3382 7814 3387
rect 6927 3339 7814 3382
rect 7808 3335 7814 3339
rect 7866 3335 7872 3387
rect 6875 3329 6927 3335
rect 3594 3318 3646 3324
rect -6846 3093 -6794 3099
rect -3972 3081 -3966 3093
rect -6794 3053 -3966 3081
rect -3972 3041 -3966 3053
rect -3914 3041 -3908 3093
rect -6846 3035 -6794 3041
rect -1792 2994 -1786 3054
rect -1726 3052 -550 3054
rect -1726 2996 -608 3052
rect -552 2996 -543 3052
rect -1726 2994 -550 2996
rect -6858 2408 -6852 2472
rect -6788 2468 -6568 2472
rect -6788 2412 -6628 2468
rect -6572 2412 -6563 2468
rect -6788 2408 -6568 2412
rect -2526 1938 -2474 1944
rect -3012 1886 -3006 1938
rect -2954 1929 -2948 1938
rect -2954 1895 -2526 1929
rect -2954 1886 -2948 1895
rect -2032 1929 -2026 1938
rect -2474 1895 -2026 1929
rect -2032 1886 -2026 1895
rect -1974 1929 -1968 1938
rect -1542 1929 -1536 1938
rect -1974 1895 -1536 1929
rect -1974 1886 -1968 1895
rect -1542 1886 -1536 1895
rect -1484 1929 -1478 1938
rect -1052 1929 -1046 1938
rect -1484 1895 -1046 1929
rect -1484 1886 -1478 1895
rect -1052 1886 -1046 1895
rect -994 1929 -988 1938
rect -532 1929 -526 1938
rect -994 1895 -526 1929
rect -994 1886 -988 1895
rect -532 1886 -526 1895
rect -474 1929 -468 1938
rect -474 1895 -443 1929
rect -474 1886 -468 1895
rect -5053 1880 -4991 1886
rect -2526 1880 -2474 1886
rect -5497 1818 -5491 1880
rect -5429 1818 -5053 1880
rect -4991 1818 -4983 1868
rect -5057 1812 -5048 1818
rect -4992 1812 -4983 1818
rect 7010 1480 7086 1489
rect 8512 1480 8588 1489
rect 7004 1416 7010 1480
rect 7086 1416 7092 1480
rect 8506 1416 8512 1480
rect 8588 1416 8594 1480
rect 7010 1407 7086 1416
rect 8512 1407 8588 1416
rect -3970 113 -3904 119
rect -5959 47 -5953 113
rect -5887 47 -3970 113
rect -3970 41 -3904 47
rect -3946 -134 -3894 -128
rect -3012 -143 -3006 -134
rect -3894 -177 -3006 -143
rect -3012 -186 -3006 -177
rect -2954 -186 -2948 -134
rect -3946 -192 -3894 -186
rect -3086 -936 -2938 -930
rect 5788 -936 5910 -930
rect -2938 -1126 -1594 -978
rect -1446 -1126 -1440 -978
rect -3086 -1174 -2938 -1168
rect 5910 -1113 7399 -991
rect 7521 -1113 7527 -991
rect 15471 -1028 15535 -1022
rect 14762 -1092 14768 -1028
rect 14832 -1092 15471 -1028
rect 15471 -1098 15535 -1092
rect 5788 -1174 5910 -1168
<< via2 >>
rect 10528 3910 10588 3914
rect 10528 3858 10532 3910
rect 10532 3858 10584 3910
rect 10584 3858 10588 3910
rect 10528 3854 10588 3858
rect -608 2996 -552 3052
rect -6628 2412 -6572 2468
rect -5048 1818 -4992 1868
rect -5048 1812 -4992 1818
rect 7010 1416 7086 1480
rect 8512 1416 8588 1480
<< metal3 >>
rect 10523 3914 10593 3919
rect 10523 3854 10528 3914
rect 10588 3854 10593 3914
rect 10523 3849 10593 3854
rect 10528 3702 10588 3849
rect -618 3638 -612 3702
rect -548 3638 -542 3702
rect 10520 3638 10526 3702
rect 10590 3638 10596 3702
rect -610 3057 -550 3638
rect -613 3052 -547 3057
rect -613 2996 -608 3052
rect -552 2996 -547 3052
rect -613 2991 -547 2996
rect 8518 2752 8582 2758
rect -5058 2688 -5052 2752
rect -4988 2688 -4982 2752
rect -6632 2592 -6568 2598
rect -6632 2473 -6568 2528
rect -6633 2468 -6567 2473
rect -6633 2412 -6628 2468
rect -6572 2412 -6567 2468
rect -6633 2407 -6567 2412
rect -5052 1873 -4988 2688
rect 7016 2592 7080 2598
rect -5053 1868 -4987 1873
rect -5053 1812 -5048 1868
rect -4992 1812 -4987 1868
rect -5053 1807 -4987 1812
rect 7016 1485 7080 2528
rect 8518 1485 8582 2688
rect 7005 1480 7091 1485
rect 7005 1416 7010 1480
rect 7086 1416 7091 1480
rect 7005 1411 7091 1416
rect 8507 1480 8593 1485
rect 8507 1416 8512 1480
rect 8588 1416 8593 1480
rect 8507 1411 8593 1416
<< via3 >>
rect -612 3638 -548 3702
rect 10526 3638 10590 3702
rect -5052 2688 -4988 2752
rect 8518 2688 8582 2752
rect -6632 2528 -6568 2592
rect 7016 2528 7080 2592
<< metal4 >>
rect -613 3702 -547 3703
rect -613 3638 -612 3702
rect -548 3700 -547 3702
rect 10525 3702 10591 3703
rect 10525 3700 10526 3702
rect -548 3640 10526 3700
rect -548 3638 -547 3640
rect -613 3637 -547 3638
rect 10525 3638 10526 3640
rect 10590 3638 10591 3702
rect 10525 3637 10591 3638
rect -5053 2752 -4987 2753
rect 8517 2752 8583 2753
rect -5053 2688 -5052 2752
rect -4988 2688 8518 2752
rect 8582 2688 8583 2752
rect -5053 2687 -4987 2688
rect 8517 2687 8583 2688
rect -6633 2592 -6567 2593
rect 7015 2592 7081 2593
rect -6633 2528 -6632 2592
rect -6568 2528 7016 2592
rect 7080 2528 7081 2592
rect -6633 2527 -6567 2528
rect 7015 2527 7081 2528
use CM_OTA_NCH  CM_OTA_NCH_0
timestamp 1710170680
transform 1 0 7260 0 1 1050
box -7100 -1050 8200 5876
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_0 ~/aicex/ip/cnr_atr_sky130nm/design/CNR_ATR_SKY130NM
timestamp 1695852000
transform 0 1 -6466 -1 0 5082
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_1
timestamp 1695852000
transform 0 1 -7456 -1 0 5082
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_2
timestamp 1695852000
transform 0 1 -6946 -1 0 5082
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_4
timestamp 1695852000
transform 0 1 -2476 -1 0 5082
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_13
timestamp 1695852000
transform 0 1 -1266 -1 0 2712
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_19
timestamp 1695852000
transform 0 1 -1756 -1 0 2712
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_20
timestamp 1695852000
transform 0 1 -5456 -1 0 5082
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_35
timestamp 1695852000
transform 0 1 -2246 -1 0 2712
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_37
timestamp 1695852000
transform 0 1 -2736 -1 0 2712
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_39
timestamp 1695852000
transform 0 1 -5976 -1 0 5082
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_41
timestamp 1695852000
transform 0 1 -746 -1 0 2712
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_59
timestamp 1695852000
transform 0 1 -3446 -1 0 5082
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_60
timestamp 1695852000
transform 0 1 -2956 -1 0 5082
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_61
timestamp 1695852000
transform 0 1 -4436 -1 0 5082
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_62
timestamp 1695852000
transform 0 1 -3936 -1 0 5082
box -184 -124 1912 613
use CNRATR_PCH_8C1F2  CNRATR_PCH_8C1F2_63
timestamp 1695852000
transform 0 1 -1476 -1 0 5092
box -184 -124 1912 613
use sky130_fd_pr__rf_pnp_05v5_W0p68L0p68  sky130_fd_pr__rf_pnp_05v5_W0p68L0p68_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1704988097
transform 1 0 -5420 0 1 800
box 0 0 796 796
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
timestamp 1704988097
transform 1 0 14840 0 1 980
box 0 0 1340 1340
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_1
timestamp 1704988097
transform 1 0 -4600 0 1 800
box 0 0 1340 1340
use SUNTR_RPPO2  SUNTR_RPPO2_1 ~/aicex/ip/cnr_gr03_sky130nm/design/SUN_TR_SKY130NM
timestamp 1710432512
transform -1 0 -2328 0 1 -4600
box 0 0 2672 4236
use SUNTR_RPPO2  SUNTR_RPPO2_2
timestamp 1710432512
transform 1 0 -7800 0 1 -4600
box 0 0 2672 4236
use SUNTR_RPPO16  SUNTR_RPPO16_0 ~/aicex/ip/cnr_gr03_sky130nm/design/SUN_TR_SKY130NM
timestamp 1710432512
transform -1 0 15520 0 1 -4600
box 0 0 8720 4236
use SUNTR_RPPO16  SUNTR_RPPO16_1
timestamp 1710432512
transform -1 0 6520 0 1 -4600
box 0 0 8720 4236
<< labels >>
flabel space -1268 4260 -1196 4324 0 FreeSans 800 0 0 0 I_OUT1
flabel metal1 -2997 -134 -2963 1886 0 FreeSans 800 0 0 0 VREF
port 2 nsew
flabel space 1180 1860 1490 1924 0 FreeSans 800 0 0 0 IBIAS
port 7 nsew
flabel locali -2245 310 17780 510 0 FreeSans 800 0 0 0 VSS
port 4 nsew
flabel locali -7412 0 18220 200 0 FreeSans 800 0 0 0 VDD
port 15 nsew
<< end >>
