*TB_SUN_TR_SKY130NM/TB_NCM
*----------------------------------------------------------------
* Include
*----------------------------------------------------------------
#ifdef Lay
.include ../../../work/lpe/TOPLEVEL_lpe.spi
#else
.include ../../../work/xsch/TOPLEVEL.spice
#endif

*-----------------------------------------------------------------
* OPTIONS
*-----------------------------------------------------------------
.option TNOM=27 GMIN=1e-15

*-----------------------------------------------------------------
* PARAMETERS
*-----------------------------------------------------------------
.param TRF = 10p

*.param AVDD = {vdda}

*-----------------------------------------------------------------
* FORCE
*-----------------------------------------------------------------
VSS  VSS  0 dc 0
VDD  VDD_1V8  VSS  dc 1.8
VRST VRST VSS PULSE(0 1.8 0.0 2NS 2NS 10US 50US)
*IBIAS VDD IBIAS dc 2u
*VRST VRST VSS dc 0


*-----------------------------------------------------------------
* DUT
*-----------------------------------------------------------------
XDUT VDD_1V8 VSS VOUT VRST TOPLEVEL

*----------------------------------------------------------------
* MEASURES
*----------------------------------------------------------------


*----------------------------------------------------------------
* PROBE
*----------------------------------------------------------------

*.save all
*TOPLEVEL valuescat
.save v(VOUT) v(VRST) v(XDUT.VREF) v(XDUT.I_PTAT) 

*Milestone 1 values
.save v(XDUT.X1.OTA_OUT) v(XDUT.X1.VD1) v(XDUT.X1.VR1)


.save i(v.XDUT.V1)
*.save all
*----------------------------------------------------------------
* NGSPICE control
*----------------------------------------------------------------
.control
set num_threads=8
set color0=white
set color1=black
unset askquit

save @m.xdut.x3.x7.xm1.msky130_fd_pr__pfet_01v8[id]

option keepopinfo
optran 0 0 0 100n 10u 0 
option keepopinfo


*ption TEMP=-40
*ran 100n 100u 30u
*rite {cicname}_-40.raw
*
*ption TEMP=0
*ran 100n 100u 30u
*rite {cicname}_0.raw

option TEMP=27
tran 10u 800u 400u


*let id = @m.xdut.x3.xm7.msky130_fd_pr__nfet_01v8[id]

write {cicname}_27.raw

*option TEMP=75
*tran 100n 100u 30u
*write {cicname}_75.raw
*
*option TEMP=125
*tran 100n 100u 30u
*write {cicname}_125.raw
*
exit

.endc

.end
