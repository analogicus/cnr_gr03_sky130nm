

.param mc_mm_switch=0
.param mc_pr_switch=0

.include tt.spi
*.include ss.spi

.lib "../../../tech/ngspice/temperature.spi" Tl

.lib "../../../tech/ngspice/supply.spi" Vl


VDD VDD 0 dc 1.8 
VSS VSS 0 dc 0


.option savecurrents
.save all
.control
optran 0 0 0 10n 10u 0
op
write MILESTONE2_TB.raw
*exit
.endc
.end
